module control_word
endmodule 