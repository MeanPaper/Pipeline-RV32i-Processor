module multiplier_control
import m_extension::*;
(
    input logic clk,
    input logic rst
);

endmodule
