// dadda_tree start here
module dadda_tree(
    input logic[31:0] opA,
    input logic[31:0] opB,
    output logic[63:0] prodAB 
);

logic [31:0] comb[32];

genvar i, j;
for(i = 0; i < 32; ++i) begin
    for(j = 0; j < 32; ++j) begin
        assign comb[i][j] = opB[i] & opA[j];
    end
end
// stage 8 begin ======================================================================================================= 
logic S_s8_280, C_s8_280;
HA HA_s8_280(.A(comb[0][28]), .B(comb[1][27]), .S(S_s8_280), .c_out(C_s8_280));
logic S_s8_290, C_s8_290;
FA FA_s8_290(.A(comb[0][29]), .B(comb[1][28]), .c_in(comb[2][27]), .S(S_s8_290), .c_out(C_s8_290));
logic S_s8_291, C_s8_291;
HA HA_s8_291(.A(comb[3][26]), .B(comb[4][25]), .S(S_s8_291), .c_out(C_s8_291));
logic S_s8_300, C_s8_300;
FA FA_s8_300(.A(comb[0][30]), .B(comb[1][29]), .c_in(comb[2][28]), .S(S_s8_300), .c_out(C_s8_300));
logic S_s8_301, C_s8_301;
FA FA_s8_301(.A(comb[3][27]), .B(comb[4][26]), .c_in(comb[5][25]), .S(S_s8_301), .c_out(C_s8_301));
logic S_s8_302, C_s8_302;
HA HA_s8_302(.A(comb[6][24]), .B(comb[7][23]), .S(S_s8_302), .c_out(C_s8_302));
logic S_s8_310, C_s8_310;
FA FA_s8_310(.A(comb[0][31]), .B(comb[1][30]), .c_in(comb[2][29]), .S(S_s8_310), .c_out(C_s8_310));
logic S_s8_311, C_s8_311;
FA FA_s8_311(.A(comb[3][28]), .B(comb[4][27]), .c_in(comb[5][26]), .S(S_s8_311), .c_out(C_s8_311));
logic S_s8_312, C_s8_312;
FA FA_s8_312(.A(comb[6][25]), .B(comb[7][24]), .c_in(comb[8][23]), .S(S_s8_312), .c_out(C_s8_312));
logic S_s8_313, C_s8_313;
HA HA_s8_313(.A(comb[9][22]), .B(comb[10][21]), .S(S_s8_313), .c_out(C_s8_313));
logic S_s8_320, C_s8_320;
FA FA_s8_320(.A(comb[1][31]), .B(comb[2][30]), .c_in(comb[3][29]), .S(S_s8_320), .c_out(C_s8_320));
logic S_s8_321, C_s8_321;
FA FA_s8_321(.A(comb[4][28]), .B(comb[5][27]), .c_in(comb[6][26]), .S(S_s8_321), .c_out(C_s8_321));
logic S_s8_322, C_s8_322;
FA FA_s8_322(.A(comb[7][25]), .B(comb[8][24]), .c_in(comb[9][23]), .S(S_s8_322), .c_out(C_s8_322));
logic S_s8_323, C_s8_323;
HA HA_s8_323(.A(comb[10][22]), .B(comb[11][21]), .S(S_s8_323), .c_out(C_s8_323));
logic S_s8_330, C_s8_330;
FA FA_s8_330(.A(comb[2][31]), .B(comb[3][30]), .c_in(comb[4][29]), .S(S_s8_330), .c_out(C_s8_330));
logic S_s8_331, C_s8_331;
FA FA_s8_331(.A(comb[5][28]), .B(comb[6][27]), .c_in(comb[7][26]), .S(S_s8_331), .c_out(C_s8_331));
logic S_s8_332, C_s8_332;
FA FA_s8_332(.A(comb[8][25]), .B(comb[9][24]), .c_in(comb[10][23]), .S(S_s8_332), .c_out(C_s8_332));
logic S_s8_340, C_s8_340;
FA FA_s8_340(.A(comb[3][31]), .B(comb[4][30]), .c_in(comb[5][29]), .S(S_s8_340), .c_out(C_s8_340));
logic S_s8_341, C_s8_341;
FA FA_s8_341(.A(comb[6][28]), .B(comb[7][27]), .c_in(comb[8][26]), .S(S_s8_341), .c_out(C_s8_341));
logic S_s8_350, C_s8_350;
FA FA_s8_350(.A(comb[4][31]), .B(comb[5][30]), .c_in(comb[6][29]), .S(S_s8_350), .c_out(C_s8_350));
// stage 8 end ======================================================================================================= 

// stage 7 begin ======================================================================================================= 
logic S_s7_190, C_s7_190;
HA HA_s7_190(.A(comb[0][19]), .B(comb[1][18]), .S(S_s7_190), .c_out(C_s7_190));
logic S_s7_200, C_s7_200;
FA FA_s7_200(.A(comb[0][20]), .B(comb[1][19]), .c_in(comb[2][18]), .S(S_s7_200), .c_out(C_s7_200));
logic S_s7_201, C_s7_201;
HA HA_s7_201(.A(comb[3][17]), .B(comb[4][16]), .S(S_s7_201), .c_out(C_s7_201));
logic S_s7_210, C_s7_210;
FA FA_s7_210(.A(comb[0][21]), .B(comb[1][20]), .c_in(comb[2][19]), .S(S_s7_210), .c_out(C_s7_210));
logic S_s7_211, C_s7_211;
FA FA_s7_211(.A(comb[3][18]), .B(comb[4][17]), .c_in(comb[5][16]), .S(S_s7_211), .c_out(C_s7_211));
logic S_s7_212, C_s7_212;
HA HA_s7_212(.A(comb[6][15]), .B(comb[7][14]), .S(S_s7_212), .c_out(C_s7_212));
logic S_s7_220, C_s7_220;
FA FA_s7_220(.A(comb[0][22]), .B(comb[1][21]), .c_in(comb[2][20]), .S(S_s7_220), .c_out(C_s7_220));
logic S_s7_221, C_s7_221;
FA FA_s7_221(.A(comb[3][19]), .B(comb[4][18]), .c_in(comb[5][17]), .S(S_s7_221), .c_out(C_s7_221));
logic S_s7_222, C_s7_222;
FA FA_s7_222(.A(comb[6][16]), .B(comb[7][15]), .c_in(comb[8][14]), .S(S_s7_222), .c_out(C_s7_222));
logic S_s7_223, C_s7_223;
HA HA_s7_223(.A(comb[9][13]), .B(comb[10][12]), .S(S_s7_223), .c_out(C_s7_223));
logic S_s7_230, C_s7_230;
FA FA_s7_230(.A(comb[0][23]), .B(comb[1][22]), .c_in(comb[2][21]), .S(S_s7_230), .c_out(C_s7_230));
logic S_s7_231, C_s7_231;
FA FA_s7_231(.A(comb[3][20]), .B(comb[4][19]), .c_in(comb[5][18]), .S(S_s7_231), .c_out(C_s7_231));
logic S_s7_232, C_s7_232;
FA FA_s7_232(.A(comb[6][17]), .B(comb[7][16]), .c_in(comb[8][15]), .S(S_s7_232), .c_out(C_s7_232));
logic S_s7_233, C_s7_233;
FA FA_s7_233(.A(comb[9][14]), .B(comb[10][13]), .c_in(comb[11][12]), .S(S_s7_233), .c_out(C_s7_233));
logic S_s7_234, C_s7_234;
HA HA_s7_234(.A(comb[12][11]), .B(comb[13][10]), .S(S_s7_234), .c_out(C_s7_234));
logic S_s7_240, C_s7_240;
FA FA_s7_240(.A(comb[0][24]), .B(comb[1][23]), .c_in(comb[2][22]), .S(S_s7_240), .c_out(C_s7_240));
logic S_s7_241, C_s7_241;
FA FA_s7_241(.A(comb[3][21]), .B(comb[4][20]), .c_in(comb[5][19]), .S(S_s7_241), .c_out(C_s7_241));
logic S_s7_242, C_s7_242;
FA FA_s7_242(.A(comb[6][18]), .B(comb[7][17]), .c_in(comb[8][16]), .S(S_s7_242), .c_out(C_s7_242));
logic S_s7_243, C_s7_243;
FA FA_s7_243(.A(comb[9][15]), .B(comb[10][14]), .c_in(comb[11][13]), .S(S_s7_243), .c_out(C_s7_243));
logic S_s7_244, C_s7_244;
FA FA_s7_244(.A(comb[12][12]), .B(comb[13][11]), .c_in(comb[14][10]), .S(S_s7_244), .c_out(C_s7_244));
logic S_s7_245, C_s7_245;
HA HA_s7_245(.A(comb[15][9]), .B(comb[16][8]), .S(S_s7_245), .c_out(C_s7_245));
logic S_s7_250, C_s7_250;
FA FA_s7_250(.A(comb[0][25]), .B(comb[1][24]), .c_in(comb[2][23]), .S(S_s7_250), .c_out(C_s7_250));
logic S_s7_251, C_s7_251;
FA FA_s7_251(.A(comb[3][22]), .B(comb[4][21]), .c_in(comb[5][20]), .S(S_s7_251), .c_out(C_s7_251));
logic S_s7_252, C_s7_252;
FA FA_s7_252(.A(comb[6][19]), .B(comb[7][18]), .c_in(comb[8][17]), .S(S_s7_252), .c_out(C_s7_252));
logic S_s7_253, C_s7_253;
FA FA_s7_253(.A(comb[9][16]), .B(comb[10][15]), .c_in(comb[11][14]), .S(S_s7_253), .c_out(C_s7_253));
logic S_s7_254, C_s7_254;
FA FA_s7_254(.A(comb[12][13]), .B(comb[13][12]), .c_in(comb[14][11]), .S(S_s7_254), .c_out(C_s7_254));
logic S_s7_255, C_s7_255;
FA FA_s7_255(.A(comb[15][10]), .B(comb[16][9]), .c_in(comb[17][8]), .S(S_s7_255), .c_out(C_s7_255));
logic S_s7_256, C_s7_256;
HA HA_s7_256(.A(comb[18][7]), .B(comb[19][6]), .S(S_s7_256), .c_out(C_s7_256));
logic S_s7_260, C_s7_260;
FA FA_s7_260(.A(comb[0][26]), .B(comb[1][25]), .c_in(comb[2][24]), .S(S_s7_260), .c_out(C_s7_260));
logic S_s7_261, C_s7_261;
FA FA_s7_261(.A(comb[3][23]), .B(comb[4][22]), .c_in(comb[5][21]), .S(S_s7_261), .c_out(C_s7_261));
logic S_s7_262, C_s7_262;
FA FA_s7_262(.A(comb[6][20]), .B(comb[7][19]), .c_in(comb[8][18]), .S(S_s7_262), .c_out(C_s7_262));
logic S_s7_263, C_s7_263;
FA FA_s7_263(.A(comb[9][17]), .B(comb[10][16]), .c_in(comb[11][15]), .S(S_s7_263), .c_out(C_s7_263));
logic S_s7_264, C_s7_264;
FA FA_s7_264(.A(comb[12][14]), .B(comb[13][13]), .c_in(comb[14][12]), .S(S_s7_264), .c_out(C_s7_264));
logic S_s7_265, C_s7_265;
FA FA_s7_265(.A(comb[15][11]), .B(comb[16][10]), .c_in(comb[17][9]), .S(S_s7_265), .c_out(C_s7_265));
logic S_s7_266, C_s7_266;
FA FA_s7_266(.A(comb[18][8]), .B(comb[19][7]), .c_in(comb[20][6]), .S(S_s7_266), .c_out(C_s7_266));
logic S_s7_267, C_s7_267;
HA HA_s7_267(.A(comb[21][5]), .B(comb[22][4]), .S(S_s7_267), .c_out(C_s7_267));
logic S_s7_270, C_s7_270;
FA FA_s7_270(.A(comb[0][27]), .B(comb[1][26]), .c_in(comb[2][25]), .S(S_s7_270), .c_out(C_s7_270));
logic S_s7_271, C_s7_271;
FA FA_s7_271(.A(comb[3][24]), .B(comb[4][23]), .c_in(comb[5][22]), .S(S_s7_271), .c_out(C_s7_271));
logic S_s7_272, C_s7_272;
FA FA_s7_272(.A(comb[6][21]), .B(comb[7][20]), .c_in(comb[8][19]), .S(S_s7_272), .c_out(C_s7_272));
logic S_s7_273, C_s7_273;
FA FA_s7_273(.A(comb[9][18]), .B(comb[10][17]), .c_in(comb[11][16]), .S(S_s7_273), .c_out(C_s7_273));
logic S_s7_274, C_s7_274;
FA FA_s7_274(.A(comb[12][15]), .B(comb[13][14]), .c_in(comb[14][13]), .S(S_s7_274), .c_out(C_s7_274));
logic S_s7_275, C_s7_275;
FA FA_s7_275(.A(comb[15][12]), .B(comb[16][11]), .c_in(comb[17][10]), .S(S_s7_275), .c_out(C_s7_275));
logic S_s7_276, C_s7_276;
FA FA_s7_276(.A(comb[18][9]), .B(comb[19][8]), .c_in(comb[20][7]), .S(S_s7_276), .c_out(C_s7_276));
logic S_s7_277, C_s7_277;
FA FA_s7_277(.A(comb[21][6]), .B(comb[22][5]), .c_in(comb[23][4]), .S(S_s7_277), .c_out(C_s7_277));
logic S_s7_278, C_s7_278;
HA HA_s7_278(.A(comb[24][3]), .B(comb[25][2]), .S(S_s7_278), .c_out(C_s7_278));
logic S_s7_280, C_s7_280;
FA FA_s7_280(.A(S_s8_280), .B(comb[2][26]), .c_in(comb[3][25]), .S(S_s7_280), .c_out(C_s7_280));
logic S_s7_281, C_s7_281;
FA FA_s7_281(.A(comb[4][24]), .B(comb[5][23]), .c_in(comb[6][22]), .S(S_s7_281), .c_out(C_s7_281));
logic S_s7_282, C_s7_282;
FA FA_s7_282(.A(comb[7][21]), .B(comb[8][20]), .c_in(comb[9][19]), .S(S_s7_282), .c_out(C_s7_282));
logic S_s7_283, C_s7_283;
FA FA_s7_283(.A(comb[10][18]), .B(comb[11][17]), .c_in(comb[12][16]), .S(S_s7_283), .c_out(C_s7_283));
logic S_s7_284, C_s7_284;
FA FA_s7_284(.A(comb[13][15]), .B(comb[14][14]), .c_in(comb[15][13]), .S(S_s7_284), .c_out(C_s7_284));
logic S_s7_285, C_s7_285;
FA FA_s7_285(.A(comb[16][12]), .B(comb[17][11]), .c_in(comb[18][10]), .S(S_s7_285), .c_out(C_s7_285));
logic S_s7_286, C_s7_286;
FA FA_s7_286(.A(comb[19][9]), .B(comb[20][8]), .c_in(comb[21][7]), .S(S_s7_286), .c_out(C_s7_286));
logic S_s7_287, C_s7_287;
FA FA_s7_287(.A(comb[22][6]), .B(comb[23][5]), .c_in(comb[24][4]), .S(S_s7_287), .c_out(C_s7_287));
logic S_s7_288, C_s7_288;
FA FA_s7_288(.A(comb[25][3]), .B(comb[26][2]), .c_in(comb[27][1]), .S(S_s7_288), .c_out(C_s7_288));
logic S_s7_290, C_s7_290;
FA FA_s7_290(.A(S_s8_291), .B(S_s8_290), .c_in(C_s8_280), .S(S_s7_290), .c_out(C_s7_290));
logic S_s7_291, C_s7_291;
FA FA_s7_291(.A(comb[5][24]), .B(comb[6][23]), .c_in(comb[7][22]), .S(S_s7_291), .c_out(C_s7_291));
logic S_s7_292, C_s7_292;
FA FA_s7_292(.A(comb[8][21]), .B(comb[9][20]), .c_in(comb[10][19]), .S(S_s7_292), .c_out(C_s7_292));
logic S_s7_293, C_s7_293;
FA FA_s7_293(.A(comb[11][18]), .B(comb[12][17]), .c_in(comb[13][16]), .S(S_s7_293), .c_out(C_s7_293));
logic S_s7_294, C_s7_294;
FA FA_s7_294(.A(comb[14][15]), .B(comb[15][14]), .c_in(comb[16][13]), .S(S_s7_294), .c_out(C_s7_294));
logic S_s7_295, C_s7_295;
FA FA_s7_295(.A(comb[17][12]), .B(comb[18][11]), .c_in(comb[19][10]), .S(S_s7_295), .c_out(C_s7_295));
logic S_s7_296, C_s7_296;
FA FA_s7_296(.A(comb[20][9]), .B(comb[21][8]), .c_in(comb[22][7]), .S(S_s7_296), .c_out(C_s7_296));
logic S_s7_297, C_s7_297;
FA FA_s7_297(.A(comb[23][6]), .B(comb[24][5]), .c_in(comb[25][4]), .S(S_s7_297), .c_out(C_s7_297));
logic S_s7_298, C_s7_298;
FA FA_s7_298(.A(comb[26][3]), .B(comb[27][2]), .c_in(comb[28][1]), .S(S_s7_298), .c_out(C_s7_298));
logic S_s7_300, C_s7_300;
FA FA_s7_300(.A(S_s8_302), .B(S_s8_301), .c_in(S_s8_300), .S(S_s7_300), .c_out(C_s7_300));
logic S_s7_301, C_s7_301;
FA FA_s7_301(.A(C_s8_291), .B(C_s8_290), .c_in(comb[8][22]), .S(S_s7_301), .c_out(C_s7_301));
logic S_s7_302, C_s7_302;
FA FA_s7_302(.A(comb[9][21]), .B(comb[10][20]), .c_in(comb[11][19]), .S(S_s7_302), .c_out(C_s7_302));
logic S_s7_303, C_s7_303;
FA FA_s7_303(.A(comb[12][18]), .B(comb[13][17]), .c_in(comb[14][16]), .S(S_s7_303), .c_out(C_s7_303));
logic S_s7_304, C_s7_304;
FA FA_s7_304(.A(comb[15][15]), .B(comb[16][14]), .c_in(comb[17][13]), .S(S_s7_304), .c_out(C_s7_304));
logic S_s7_305, C_s7_305;
FA FA_s7_305(.A(comb[18][12]), .B(comb[19][11]), .c_in(comb[20][10]), .S(S_s7_305), .c_out(C_s7_305));
logic S_s7_306, C_s7_306;
FA FA_s7_306(.A(comb[21][9]), .B(comb[22][8]), .c_in(comb[23][7]), .S(S_s7_306), .c_out(C_s7_306));
logic S_s7_307, C_s7_307;
FA FA_s7_307(.A(comb[24][6]), .B(comb[25][5]), .c_in(comb[26][4]), .S(S_s7_307), .c_out(C_s7_307));
logic S_s7_308, C_s7_308;
FA FA_s7_308(.A(comb[27][3]), .B(comb[28][2]), .c_in(comb[29][1]), .S(S_s7_308), .c_out(C_s7_308));
logic S_s7_310, C_s7_310;
FA FA_s7_310(.A(S_s8_313), .B(S_s8_312), .c_in(S_s8_311), .S(S_s7_310), .c_out(C_s7_310));
logic S_s7_311, C_s7_311;
FA FA_s7_311(.A(S_s8_310), .B(C_s8_302), .c_in(C_s8_301), .S(S_s7_311), .c_out(C_s7_311));
logic S_s7_312, C_s7_312;
FA FA_s7_312(.A(C_s8_300), .B(comb[11][20]), .c_in(comb[12][19]), .S(S_s7_312), .c_out(C_s7_312));
logic S_s7_313, C_s7_313;
FA FA_s7_313(.A(comb[13][18]), .B(comb[14][17]), .c_in(comb[15][16]), .S(S_s7_313), .c_out(C_s7_313));
logic S_s7_314, C_s7_314;
FA FA_s7_314(.A(comb[16][15]), .B(comb[17][14]), .c_in(comb[18][13]), .S(S_s7_314), .c_out(C_s7_314));
logic S_s7_315, C_s7_315;
FA FA_s7_315(.A(comb[19][12]), .B(comb[20][11]), .c_in(comb[21][10]), .S(S_s7_315), .c_out(C_s7_315));
logic S_s7_316, C_s7_316;
FA FA_s7_316(.A(comb[22][9]), .B(comb[23][8]), .c_in(comb[24][7]), .S(S_s7_316), .c_out(C_s7_316));
logic S_s7_317, C_s7_317;
FA FA_s7_317(.A(comb[25][6]), .B(comb[26][5]), .c_in(comb[27][4]), .S(S_s7_317), .c_out(C_s7_317));
logic S_s7_318, C_s7_318;
FA FA_s7_318(.A(comb[28][3]), .B(comb[29][2]), .c_in(comb[30][1]), .S(S_s7_318), .c_out(C_s7_318));
logic S_s7_320, C_s7_320;
FA FA_s7_320(.A(S_s8_323), .B(S_s8_322), .c_in(S_s8_321), .S(S_s7_320), .c_out(C_s7_320));
logic S_s7_321, C_s7_321;
FA FA_s7_321(.A(S_s8_320), .B(C_s8_313), .c_in(C_s8_312), .S(S_s7_321), .c_out(C_s7_321));
logic S_s7_322, C_s7_322;
FA FA_s7_322(.A(C_s8_311), .B(C_s8_310), .c_in(comb[12][20]), .S(S_s7_322), .c_out(C_s7_322));
logic S_s7_323, C_s7_323;
FA FA_s7_323(.A(comb[13][19]), .B(comb[14][18]), .c_in(comb[15][17]), .S(S_s7_323), .c_out(C_s7_323));
logic S_s7_324, C_s7_324;
FA FA_s7_324(.A(comb[16][16]), .B(comb[17][15]), .c_in(comb[18][14]), .S(S_s7_324), .c_out(C_s7_324));
logic S_s7_325, C_s7_325;
FA FA_s7_325(.A(comb[19][13]), .B(comb[20][12]), .c_in(comb[21][11]), .S(S_s7_325), .c_out(C_s7_325));
logic S_s7_326, C_s7_326;
FA FA_s7_326(.A(comb[22][10]), .B(comb[23][9]), .c_in(comb[24][8]), .S(S_s7_326), .c_out(C_s7_326));
logic S_s7_327, C_s7_327;
FA FA_s7_327(.A(comb[25][7]), .B(comb[26][6]), .c_in(comb[27][5]), .S(S_s7_327), .c_out(C_s7_327));
logic S_s7_328, C_s7_328;
FA FA_s7_328(.A(comb[28][4]), .B(comb[29][3]), .c_in(comb[30][2]), .S(S_s7_328), .c_out(C_s7_328));
logic S_s7_330, C_s7_330;
FA FA_s7_330(.A(S_s8_332), .B(S_s8_331), .c_in(S_s8_330), .S(S_s7_330), .c_out(C_s7_330));
logic S_s7_331, C_s7_331;
FA FA_s7_331(.A(C_s8_323), .B(C_s8_322), .c_in(C_s8_321), .S(S_s7_331), .c_out(C_s7_331));
logic S_s7_332, C_s7_332;
FA FA_s7_332(.A(C_s8_320), .B(comb[11][22]), .c_in(comb[12][21]), .S(S_s7_332), .c_out(C_s7_332));
logic S_s7_333, C_s7_333;
FA FA_s7_333(.A(comb[13][20]), .B(comb[14][19]), .c_in(comb[15][18]), .S(S_s7_333), .c_out(C_s7_333));
logic S_s7_334, C_s7_334;
FA FA_s7_334(.A(comb[16][17]), .B(comb[17][16]), .c_in(comb[18][15]), .S(S_s7_334), .c_out(C_s7_334));
logic S_s7_335, C_s7_335;
FA FA_s7_335(.A(comb[19][14]), .B(comb[20][13]), .c_in(comb[21][12]), .S(S_s7_335), .c_out(C_s7_335));
logic S_s7_336, C_s7_336;
FA FA_s7_336(.A(comb[22][11]), .B(comb[23][10]), .c_in(comb[24][9]), .S(S_s7_336), .c_out(C_s7_336));
logic S_s7_337, C_s7_337;
FA FA_s7_337(.A(comb[25][8]), .B(comb[26][7]), .c_in(comb[27][6]), .S(S_s7_337), .c_out(C_s7_337));
logic S_s7_338, C_s7_338;
FA FA_s7_338(.A(comb[28][5]), .B(comb[29][4]), .c_in(comb[30][3]), .S(S_s7_338), .c_out(C_s7_338));
logic S_s7_340, C_s7_340;
FA FA_s7_340(.A(S_s8_341), .B(S_s8_340), .c_in(C_s8_332), .S(S_s7_340), .c_out(C_s7_340));
logic S_s7_341, C_s7_341;
FA FA_s7_341(.A(C_s8_331), .B(C_s8_330), .c_in(comb[9][25]), .S(S_s7_341), .c_out(C_s7_341));
logic S_s7_342, C_s7_342;
FA FA_s7_342(.A(comb[10][24]), .B(comb[11][23]), .c_in(comb[12][22]), .S(S_s7_342), .c_out(C_s7_342));
logic S_s7_343, C_s7_343;
FA FA_s7_343(.A(comb[13][21]), .B(comb[14][20]), .c_in(comb[15][19]), .S(S_s7_343), .c_out(C_s7_343));
logic S_s7_344, C_s7_344;
FA FA_s7_344(.A(comb[16][18]), .B(comb[17][17]), .c_in(comb[18][16]), .S(S_s7_344), .c_out(C_s7_344));
logic S_s7_345, C_s7_345;
FA FA_s7_345(.A(comb[19][15]), .B(comb[20][14]), .c_in(comb[21][13]), .S(S_s7_345), .c_out(C_s7_345));
logic S_s7_346, C_s7_346;
FA FA_s7_346(.A(comb[22][12]), .B(comb[23][11]), .c_in(comb[24][10]), .S(S_s7_346), .c_out(C_s7_346));
logic S_s7_347, C_s7_347;
FA FA_s7_347(.A(comb[25][9]), .B(comb[26][8]), .c_in(comb[27][7]), .S(S_s7_347), .c_out(C_s7_347));
logic S_s7_348, C_s7_348;
FA FA_s7_348(.A(comb[28][6]), .B(comb[29][5]), .c_in(comb[30][4]), .S(S_s7_348), .c_out(C_s7_348));
logic S_s7_350, C_s7_350;
FA FA_s7_350(.A(S_s8_350), .B(C_s8_341), .c_in(C_s8_340), .S(S_s7_350), .c_out(C_s7_350));
logic S_s7_351, C_s7_351;
FA FA_s7_351(.A(comb[7][28]), .B(comb[8][27]), .c_in(comb[9][26]), .S(S_s7_351), .c_out(C_s7_351));
logic S_s7_352, C_s7_352;
FA FA_s7_352(.A(comb[10][25]), .B(comb[11][24]), .c_in(comb[12][23]), .S(S_s7_352), .c_out(C_s7_352));
logic S_s7_353, C_s7_353;
FA FA_s7_353(.A(comb[13][22]), .B(comb[14][21]), .c_in(comb[15][20]), .S(S_s7_353), .c_out(C_s7_353));
logic S_s7_354, C_s7_354;
FA FA_s7_354(.A(comb[16][19]), .B(comb[17][18]), .c_in(comb[18][17]), .S(S_s7_354), .c_out(C_s7_354));
logic S_s7_355, C_s7_355;
FA FA_s7_355(.A(comb[19][16]), .B(comb[20][15]), .c_in(comb[21][14]), .S(S_s7_355), .c_out(C_s7_355));
logic S_s7_356, C_s7_356;
FA FA_s7_356(.A(comb[22][13]), .B(comb[23][12]), .c_in(comb[24][11]), .S(S_s7_356), .c_out(C_s7_356));
logic S_s7_357, C_s7_357;
FA FA_s7_357(.A(comb[25][10]), .B(comb[26][9]), .c_in(comb[27][8]), .S(S_s7_357), .c_out(C_s7_357));
logic S_s7_358, C_s7_358;
FA FA_s7_358(.A(comb[28][7]), .B(comb[29][6]), .c_in(comb[30][5]), .S(S_s7_358), .c_out(C_s7_358));
logic S_s7_360, C_s7_360;
FA FA_s7_360(.A(C_s8_350), .B(comb[5][31]), .c_in(comb[6][30]), .S(S_s7_360), .c_out(C_s7_360));
logic S_s7_361, C_s7_361;
FA FA_s7_361(.A(comb[7][29]), .B(comb[8][28]), .c_in(comb[9][27]), .S(S_s7_361), .c_out(C_s7_361));
logic S_s7_362, C_s7_362;
FA FA_s7_362(.A(comb[10][26]), .B(comb[11][25]), .c_in(comb[12][24]), .S(S_s7_362), .c_out(C_s7_362));
logic S_s7_363, C_s7_363;
FA FA_s7_363(.A(comb[13][23]), .B(comb[14][22]), .c_in(comb[15][21]), .S(S_s7_363), .c_out(C_s7_363));
logic S_s7_364, C_s7_364;
FA FA_s7_364(.A(comb[16][20]), .B(comb[17][19]), .c_in(comb[18][18]), .S(S_s7_364), .c_out(C_s7_364));
logic S_s7_365, C_s7_365;
FA FA_s7_365(.A(comb[19][17]), .B(comb[20][16]), .c_in(comb[21][15]), .S(S_s7_365), .c_out(C_s7_365));
logic S_s7_366, C_s7_366;
FA FA_s7_366(.A(comb[22][14]), .B(comb[23][13]), .c_in(comb[24][12]), .S(S_s7_366), .c_out(C_s7_366));
logic S_s7_367, C_s7_367;
FA FA_s7_367(.A(comb[25][11]), .B(comb[26][10]), .c_in(comb[27][9]), .S(S_s7_367), .c_out(C_s7_367));
logic S_s7_368, C_s7_368;
FA FA_s7_368(.A(comb[28][8]), .B(comb[29][7]), .c_in(comb[30][6]), .S(S_s7_368), .c_out(C_s7_368));
logic S_s7_370, C_s7_370;
FA FA_s7_370(.A(comb[6][31]), .B(comb[7][30]), .c_in(comb[8][29]), .S(S_s7_370), .c_out(C_s7_370));
logic S_s7_371, C_s7_371;
FA FA_s7_371(.A(comb[9][28]), .B(comb[10][27]), .c_in(comb[11][26]), .S(S_s7_371), .c_out(C_s7_371));
logic S_s7_372, C_s7_372;
FA FA_s7_372(.A(comb[12][25]), .B(comb[13][24]), .c_in(comb[14][23]), .S(S_s7_372), .c_out(C_s7_372));
logic S_s7_373, C_s7_373;
FA FA_s7_373(.A(comb[15][22]), .B(comb[16][21]), .c_in(comb[17][20]), .S(S_s7_373), .c_out(C_s7_373));
logic S_s7_374, C_s7_374;
FA FA_s7_374(.A(comb[18][19]), .B(comb[19][18]), .c_in(comb[20][17]), .S(S_s7_374), .c_out(C_s7_374));
logic S_s7_375, C_s7_375;
FA FA_s7_375(.A(comb[21][16]), .B(comb[22][15]), .c_in(comb[23][14]), .S(S_s7_375), .c_out(C_s7_375));
logic S_s7_376, C_s7_376;
FA FA_s7_376(.A(comb[24][13]), .B(comb[25][12]), .c_in(comb[26][11]), .S(S_s7_376), .c_out(C_s7_376));
logic S_s7_377, C_s7_377;
FA FA_s7_377(.A(comb[27][10]), .B(comb[28][9]), .c_in(comb[29][8]), .S(S_s7_377), .c_out(C_s7_377));
logic S_s7_380, C_s7_380;
FA FA_s7_380(.A(comb[7][31]), .B(comb[8][30]), .c_in(comb[9][29]), .S(S_s7_380), .c_out(C_s7_380));
logic S_s7_381, C_s7_381;
FA FA_s7_381(.A(comb[10][28]), .B(comb[11][27]), .c_in(comb[12][26]), .S(S_s7_381), .c_out(C_s7_381));
logic S_s7_382, C_s7_382;
FA FA_s7_382(.A(comb[13][25]), .B(comb[14][24]), .c_in(comb[15][23]), .S(S_s7_382), .c_out(C_s7_382));
logic S_s7_383, C_s7_383;
FA FA_s7_383(.A(comb[16][22]), .B(comb[17][21]), .c_in(comb[18][20]), .S(S_s7_383), .c_out(C_s7_383));
logic S_s7_384, C_s7_384;
FA FA_s7_384(.A(comb[19][19]), .B(comb[20][18]), .c_in(comb[21][17]), .S(S_s7_384), .c_out(C_s7_384));
logic S_s7_385, C_s7_385;
FA FA_s7_385(.A(comb[22][16]), .B(comb[23][15]), .c_in(comb[24][14]), .S(S_s7_385), .c_out(C_s7_385));
logic S_s7_386, C_s7_386;
FA FA_s7_386(.A(comb[25][13]), .B(comb[26][12]), .c_in(comb[27][11]), .S(S_s7_386), .c_out(C_s7_386));
logic S_s7_390, C_s7_390;
FA FA_s7_390(.A(comb[8][31]), .B(comb[9][30]), .c_in(comb[10][29]), .S(S_s7_390), .c_out(C_s7_390));
logic S_s7_391, C_s7_391;
FA FA_s7_391(.A(comb[11][28]), .B(comb[12][27]), .c_in(comb[13][26]), .S(S_s7_391), .c_out(C_s7_391));
logic S_s7_392, C_s7_392;
FA FA_s7_392(.A(comb[14][25]), .B(comb[15][24]), .c_in(comb[16][23]), .S(S_s7_392), .c_out(C_s7_392));
logic S_s7_393, C_s7_393;
FA FA_s7_393(.A(comb[17][22]), .B(comb[18][21]), .c_in(comb[19][20]), .S(S_s7_393), .c_out(C_s7_393));
logic S_s7_394, C_s7_394;
FA FA_s7_394(.A(comb[20][19]), .B(comb[21][18]), .c_in(comb[22][17]), .S(S_s7_394), .c_out(C_s7_394));
logic S_s7_395, C_s7_395;
FA FA_s7_395(.A(comb[23][16]), .B(comb[24][15]), .c_in(comb[25][14]), .S(S_s7_395), .c_out(C_s7_395));
logic S_s7_400, C_s7_400;
FA FA_s7_400(.A(comb[9][31]), .B(comb[10][30]), .c_in(comb[11][29]), .S(S_s7_400), .c_out(C_s7_400));
logic S_s7_401, C_s7_401;
FA FA_s7_401(.A(comb[12][28]), .B(comb[13][27]), .c_in(comb[14][26]), .S(S_s7_401), .c_out(C_s7_401));
logic S_s7_402, C_s7_402;
FA FA_s7_402(.A(comb[15][25]), .B(comb[16][24]), .c_in(comb[17][23]), .S(S_s7_402), .c_out(C_s7_402));
logic S_s7_403, C_s7_403;
FA FA_s7_403(.A(comb[18][22]), .B(comb[19][21]), .c_in(comb[20][20]), .S(S_s7_403), .c_out(C_s7_403));
logic S_s7_404, C_s7_404;
FA FA_s7_404(.A(comb[21][19]), .B(comb[22][18]), .c_in(comb[23][17]), .S(S_s7_404), .c_out(C_s7_404));
logic S_s7_410, C_s7_410;
FA FA_s7_410(.A(comb[10][31]), .B(comb[11][30]), .c_in(comb[12][29]), .S(S_s7_410), .c_out(C_s7_410));
logic S_s7_411, C_s7_411;
FA FA_s7_411(.A(comb[13][28]), .B(comb[14][27]), .c_in(comb[15][26]), .S(S_s7_411), .c_out(C_s7_411));
logic S_s7_412, C_s7_412;
FA FA_s7_412(.A(comb[16][25]), .B(comb[17][24]), .c_in(comb[18][23]), .S(S_s7_412), .c_out(C_s7_412));
logic S_s7_413, C_s7_413;
FA FA_s7_413(.A(comb[19][22]), .B(comb[20][21]), .c_in(comb[21][20]), .S(S_s7_413), .c_out(C_s7_413));
logic S_s7_420, C_s7_420;
FA FA_s7_420(.A(comb[11][31]), .B(comb[12][30]), .c_in(comb[13][29]), .S(S_s7_420), .c_out(C_s7_420));
logic S_s7_421, C_s7_421;
FA FA_s7_421(.A(comb[14][28]), .B(comb[15][27]), .c_in(comb[16][26]), .S(S_s7_421), .c_out(C_s7_421));
logic S_s7_422, C_s7_422;
FA FA_s7_422(.A(comb[17][25]), .B(comb[18][24]), .c_in(comb[19][23]), .S(S_s7_422), .c_out(C_s7_422));
logic S_s7_430, C_s7_430;
FA FA_s7_430(.A(comb[12][31]), .B(comb[13][30]), .c_in(comb[14][29]), .S(S_s7_430), .c_out(C_s7_430));
logic S_s7_431, C_s7_431;
FA FA_s7_431(.A(comb[15][28]), .B(comb[16][27]), .c_in(comb[17][26]), .S(S_s7_431), .c_out(C_s7_431));
logic S_s7_440, C_s7_440;
FA FA_s7_440(.A(comb[13][31]), .B(comb[14][30]), .c_in(comb[15][29]), .S(S_s7_440), .c_out(C_s7_440));
// stage 7 end ======================================================================================================= 

// stage 6 begin ======================================================================================================= 
logic S_s6_130, C_s6_130;
HA HA_s6_130(.A(comb[0][13]), .B(comb[1][12]), .S(S_s6_130), .c_out(C_s6_130));
logic S_s6_140, C_s6_140;
FA FA_s6_140(.A(comb[0][14]), .B(comb[1][13]), .c_in(comb[2][12]), .S(S_s6_140), .c_out(C_s6_140));
logic S_s6_141, C_s6_141;
HA HA_s6_141(.A(comb[3][11]), .B(comb[4][10]), .S(S_s6_141), .c_out(C_s6_141));
logic S_s6_150, C_s6_150;
FA FA_s6_150(.A(comb[0][15]), .B(comb[1][14]), .c_in(comb[2][13]), .S(S_s6_150), .c_out(C_s6_150));
logic S_s6_151, C_s6_151;
FA FA_s6_151(.A(comb[3][12]), .B(comb[4][11]), .c_in(comb[5][10]), .S(S_s6_151), .c_out(C_s6_151));
logic S_s6_152, C_s6_152;
HA HA_s6_152(.A(comb[6][9]), .B(comb[7][8]), .S(S_s6_152), .c_out(C_s6_152));
logic S_s6_160, C_s6_160;
FA FA_s6_160(.A(comb[0][16]), .B(comb[1][15]), .c_in(comb[2][14]), .S(S_s6_160), .c_out(C_s6_160));
logic S_s6_161, C_s6_161;
FA FA_s6_161(.A(comb[3][13]), .B(comb[4][12]), .c_in(comb[5][11]), .S(S_s6_161), .c_out(C_s6_161));
logic S_s6_162, C_s6_162;
FA FA_s6_162(.A(comb[6][10]), .B(comb[7][9]), .c_in(comb[8][8]), .S(S_s6_162), .c_out(C_s6_162));
logic S_s6_163, C_s6_163;
HA HA_s6_163(.A(comb[9][7]), .B(comb[10][6]), .S(S_s6_163), .c_out(C_s6_163));
logic S_s6_170, C_s6_170;
FA FA_s6_170(.A(comb[0][17]), .B(comb[1][16]), .c_in(comb[2][15]), .S(S_s6_170), .c_out(C_s6_170));
logic S_s6_171, C_s6_171;
FA FA_s6_171(.A(comb[3][14]), .B(comb[4][13]), .c_in(comb[5][12]), .S(S_s6_171), .c_out(C_s6_171));
logic S_s6_172, C_s6_172;
FA FA_s6_172(.A(comb[6][11]), .B(comb[7][10]), .c_in(comb[8][9]), .S(S_s6_172), .c_out(C_s6_172));
logic S_s6_173, C_s6_173;
FA FA_s6_173(.A(comb[9][8]), .B(comb[10][7]), .c_in(comb[11][6]), .S(S_s6_173), .c_out(C_s6_173));
logic S_s6_174, C_s6_174;
HA HA_s6_174(.A(comb[12][5]), .B(comb[13][4]), .S(S_s6_174), .c_out(C_s6_174));
logic S_s6_180, C_s6_180;
FA FA_s6_180(.A(comb[0][18]), .B(comb[1][17]), .c_in(comb[2][16]), .S(S_s6_180), .c_out(C_s6_180));
logic S_s6_181, C_s6_181;
FA FA_s6_181(.A(comb[3][15]), .B(comb[4][14]), .c_in(comb[5][13]), .S(S_s6_181), .c_out(C_s6_181));
logic S_s6_182, C_s6_182;
FA FA_s6_182(.A(comb[6][12]), .B(comb[7][11]), .c_in(comb[8][10]), .S(S_s6_182), .c_out(C_s6_182));
logic S_s6_183, C_s6_183;
FA FA_s6_183(.A(comb[9][9]), .B(comb[10][8]), .c_in(comb[11][7]), .S(S_s6_183), .c_out(C_s6_183));
logic S_s6_184, C_s6_184;
FA FA_s6_184(.A(comb[12][6]), .B(comb[13][5]), .c_in(comb[14][4]), .S(S_s6_184), .c_out(C_s6_184));
logic S_s6_185, C_s6_185;
HA HA_s6_185(.A(comb[15][3]), .B(comb[16][2]), .S(S_s6_185), .c_out(C_s6_185));
logic S_s6_190, C_s6_190;
FA FA_s6_190(.A(S_s7_190), .B(comb[2][17]), .c_in(comb[3][16]), .S(S_s6_190), .c_out(C_s6_190));
logic S_s6_191, C_s6_191;
FA FA_s6_191(.A(comb[4][15]), .B(comb[5][14]), .c_in(comb[6][13]), .S(S_s6_191), .c_out(C_s6_191));
logic S_s6_192, C_s6_192;
FA FA_s6_192(.A(comb[7][12]), .B(comb[8][11]), .c_in(comb[9][10]), .S(S_s6_192), .c_out(C_s6_192));
logic S_s6_193, C_s6_193;
FA FA_s6_193(.A(comb[10][9]), .B(comb[11][8]), .c_in(comb[12][7]), .S(S_s6_193), .c_out(C_s6_193));
logic S_s6_194, C_s6_194;
FA FA_s6_194(.A(comb[13][6]), .B(comb[14][5]), .c_in(comb[15][4]), .S(S_s6_194), .c_out(C_s6_194));
logic S_s6_195, C_s6_195;
FA FA_s6_195(.A(comb[16][3]), .B(comb[17][2]), .c_in(comb[18][1]), .S(S_s6_195), .c_out(C_s6_195));
logic S_s6_200, C_s6_200;
FA FA_s6_200(.A(S_s7_201), .B(S_s7_200), .c_in(C_s7_190), .S(S_s6_200), .c_out(C_s6_200));
logic S_s6_201, C_s6_201;
FA FA_s6_201(.A(comb[5][15]), .B(comb[6][14]), .c_in(comb[7][13]), .S(S_s6_201), .c_out(C_s6_201));
logic S_s6_202, C_s6_202;
FA FA_s6_202(.A(comb[8][12]), .B(comb[9][11]), .c_in(comb[10][10]), .S(S_s6_202), .c_out(C_s6_202));
logic S_s6_203, C_s6_203;
FA FA_s6_203(.A(comb[11][9]), .B(comb[12][8]), .c_in(comb[13][7]), .S(S_s6_203), .c_out(C_s6_203));
logic S_s6_204, C_s6_204;
FA FA_s6_204(.A(comb[14][6]), .B(comb[15][5]), .c_in(comb[16][4]), .S(S_s6_204), .c_out(C_s6_204));
logic S_s6_205, C_s6_205;
FA FA_s6_205(.A(comb[17][3]), .B(comb[18][2]), .c_in(comb[19][1]), .S(S_s6_205), .c_out(C_s6_205));
logic S_s6_210, C_s6_210;
FA FA_s6_210(.A(S_s7_212), .B(S_s7_211), .c_in(S_s7_210), .S(S_s6_210), .c_out(C_s6_210));
logic S_s6_211, C_s6_211;
FA FA_s6_211(.A(C_s7_201), .B(C_s7_200), .c_in(comb[8][13]), .S(S_s6_211), .c_out(C_s6_211));
logic S_s6_212, C_s6_212;
FA FA_s6_212(.A(comb[9][12]), .B(comb[10][11]), .c_in(comb[11][10]), .S(S_s6_212), .c_out(C_s6_212));
logic S_s6_213, C_s6_213;
FA FA_s6_213(.A(comb[12][9]), .B(comb[13][8]), .c_in(comb[14][7]), .S(S_s6_213), .c_out(C_s6_213));
logic S_s6_214, C_s6_214;
FA FA_s6_214(.A(comb[15][6]), .B(comb[16][5]), .c_in(comb[17][4]), .S(S_s6_214), .c_out(C_s6_214));
logic S_s6_215, C_s6_215;
FA FA_s6_215(.A(comb[18][3]), .B(comb[19][2]), .c_in(comb[20][1]), .S(S_s6_215), .c_out(C_s6_215));
logic S_s6_220, C_s6_220;
FA FA_s6_220(.A(S_s7_223), .B(S_s7_222), .c_in(S_s7_221), .S(S_s6_220), .c_out(C_s6_220));
logic S_s6_221, C_s6_221;
FA FA_s6_221(.A(S_s7_220), .B(C_s7_212), .c_in(C_s7_211), .S(S_s6_221), .c_out(C_s6_221));
logic S_s6_222, C_s6_222;
FA FA_s6_222(.A(C_s7_210), .B(comb[11][11]), .c_in(comb[12][10]), .S(S_s6_222), .c_out(C_s6_222));
logic S_s6_223, C_s6_223;
FA FA_s6_223(.A(comb[13][9]), .B(comb[14][8]), .c_in(comb[15][7]), .S(S_s6_223), .c_out(C_s6_223));
logic S_s6_224, C_s6_224;
FA FA_s6_224(.A(comb[16][6]), .B(comb[17][5]), .c_in(comb[18][4]), .S(S_s6_224), .c_out(C_s6_224));
logic S_s6_225, C_s6_225;
FA FA_s6_225(.A(comb[19][3]), .B(comb[20][2]), .c_in(comb[21][1]), .S(S_s6_225), .c_out(C_s6_225));
logic S_s6_230, C_s6_230;
FA FA_s6_230(.A(S_s7_234), .B(S_s7_233), .c_in(S_s7_232), .S(S_s6_230), .c_out(C_s6_230));
logic S_s6_231, C_s6_231;
FA FA_s6_231(.A(S_s7_231), .B(S_s7_230), .c_in(C_s7_223), .S(S_s6_231), .c_out(C_s6_231));
logic S_s6_232, C_s6_232;
FA FA_s6_232(.A(C_s7_222), .B(C_s7_221), .c_in(C_s7_220), .S(S_s6_232), .c_out(C_s6_232));
logic S_s6_233, C_s6_233;
FA FA_s6_233(.A(comb[14][9]), .B(comb[15][8]), .c_in(comb[16][7]), .S(S_s6_233), .c_out(C_s6_233));
logic S_s6_234, C_s6_234;
FA FA_s6_234(.A(comb[17][6]), .B(comb[18][5]), .c_in(comb[19][4]), .S(S_s6_234), .c_out(C_s6_234));
logic S_s6_235, C_s6_235;
FA FA_s6_235(.A(comb[20][3]), .B(comb[21][2]), .c_in(comb[22][1]), .S(S_s6_235), .c_out(C_s6_235));
logic S_s6_240, C_s6_240;
FA FA_s6_240(.A(S_s7_245), .B(S_s7_244), .c_in(S_s7_243), .S(S_s6_240), .c_out(C_s6_240));
logic S_s6_241, C_s6_241;
FA FA_s6_241(.A(S_s7_242), .B(S_s7_241), .c_in(S_s7_240), .S(S_s6_241), .c_out(C_s6_241));
logic S_s6_242, C_s6_242;
FA FA_s6_242(.A(C_s7_234), .B(C_s7_233), .c_in(C_s7_232), .S(S_s6_242), .c_out(C_s6_242));
logic S_s6_243, C_s6_243;
FA FA_s6_243(.A(C_s7_231), .B(C_s7_230), .c_in(comb[17][7]), .S(S_s6_243), .c_out(C_s6_243));
logic S_s6_244, C_s6_244;
FA FA_s6_244(.A(comb[18][6]), .B(comb[19][5]), .c_in(comb[20][4]), .S(S_s6_244), .c_out(C_s6_244));
logic S_s6_245, C_s6_245;
FA FA_s6_245(.A(comb[21][3]), .B(comb[22][2]), .c_in(comb[23][1]), .S(S_s6_245), .c_out(C_s6_245));
logic S_s6_250, C_s6_250;
FA FA_s6_250(.A(S_s7_256), .B(S_s7_255), .c_in(S_s7_254), .S(S_s6_250), .c_out(C_s6_250));
logic S_s6_251, C_s6_251;
FA FA_s6_251(.A(S_s7_253), .B(S_s7_252), .c_in(S_s7_251), .S(S_s6_251), .c_out(C_s6_251));
logic S_s6_252, C_s6_252;
FA FA_s6_252(.A(S_s7_250), .B(C_s7_245), .c_in(C_s7_244), .S(S_s6_252), .c_out(C_s6_252));
logic S_s6_253, C_s6_253;
FA FA_s6_253(.A(C_s7_243), .B(C_s7_242), .c_in(C_s7_241), .S(S_s6_253), .c_out(C_s6_253));
logic S_s6_254, C_s6_254;
FA FA_s6_254(.A(C_s7_240), .B(comb[20][5]), .c_in(comb[21][4]), .S(S_s6_254), .c_out(C_s6_254));
logic S_s6_255, C_s6_255;
FA FA_s6_255(.A(comb[22][3]), .B(comb[23][2]), .c_in(comb[24][1]), .S(S_s6_255), .c_out(C_s6_255));
logic S_s6_260, C_s6_260;
FA FA_s6_260(.A(S_s7_267), .B(S_s7_266), .c_in(S_s7_265), .S(S_s6_260), .c_out(C_s6_260));
logic S_s6_261, C_s6_261;
FA FA_s6_261(.A(S_s7_264), .B(S_s7_263), .c_in(S_s7_262), .S(S_s6_261), .c_out(C_s6_261));
logic S_s6_262, C_s6_262;
FA FA_s6_262(.A(S_s7_261), .B(S_s7_260), .c_in(C_s7_256), .S(S_s6_262), .c_out(C_s6_262));
logic S_s6_263, C_s6_263;
FA FA_s6_263(.A(C_s7_255), .B(C_s7_254), .c_in(C_s7_253), .S(S_s6_263), .c_out(C_s6_263));
logic S_s6_264, C_s6_264;
FA FA_s6_264(.A(C_s7_252), .B(C_s7_251), .c_in(C_s7_250), .S(S_s6_264), .c_out(C_s6_264));
logic S_s6_265, C_s6_265;
FA FA_s6_265(.A(comb[23][3]), .B(comb[24][2]), .c_in(comb[25][1]), .S(S_s6_265), .c_out(C_s6_265));
logic S_s6_270, C_s6_270;
FA FA_s6_270(.A(S_s7_278), .B(S_s7_277), .c_in(S_s7_276), .S(S_s6_270), .c_out(C_s6_270));
logic S_s6_271, C_s6_271;
FA FA_s6_271(.A(S_s7_275), .B(S_s7_274), .c_in(S_s7_273), .S(S_s6_271), .c_out(C_s6_271));
logic S_s6_272, C_s6_272;
FA FA_s6_272(.A(S_s7_272), .B(S_s7_271), .c_in(S_s7_270), .S(S_s6_272), .c_out(C_s6_272));
logic S_s6_273, C_s6_273;
FA FA_s6_273(.A(C_s7_267), .B(C_s7_266), .c_in(C_s7_265), .S(S_s6_273), .c_out(C_s6_273));
logic S_s6_274, C_s6_274;
FA FA_s6_274(.A(C_s7_264), .B(C_s7_263), .c_in(C_s7_262), .S(S_s6_274), .c_out(C_s6_274));
logic S_s6_275, C_s6_275;
FA FA_s6_275(.A(C_s7_261), .B(C_s7_260), .c_in(comb[26][1]), .S(S_s6_275), .c_out(C_s6_275));
logic S_s6_280, C_s6_280;
FA FA_s6_280(.A(S_s7_288), .B(S_s7_287), .c_in(S_s7_286), .S(S_s6_280), .c_out(C_s6_280));
logic S_s6_281, C_s6_281;
FA FA_s6_281(.A(S_s7_285), .B(S_s7_284), .c_in(S_s7_283), .S(S_s6_281), .c_out(C_s6_281));
logic S_s6_282, C_s6_282;
FA FA_s6_282(.A(S_s7_282), .B(S_s7_281), .c_in(S_s7_280), .S(S_s6_282), .c_out(C_s6_282));
logic S_s6_283, C_s6_283;
FA FA_s6_283(.A(C_s7_278), .B(C_s7_277), .c_in(C_s7_276), .S(S_s6_283), .c_out(C_s6_283));
logic S_s6_284, C_s6_284;
FA FA_s6_284(.A(C_s7_275), .B(C_s7_274), .c_in(C_s7_273), .S(S_s6_284), .c_out(C_s6_284));
logic S_s6_285, C_s6_285;
FA FA_s6_285(.A(C_s7_272), .B(C_s7_271), .c_in(C_s7_270), .S(S_s6_285), .c_out(C_s6_285));
logic S_s6_290, C_s6_290;
FA FA_s6_290(.A(S_s7_298), .B(S_s7_297), .c_in(S_s7_296), .S(S_s6_290), .c_out(C_s6_290));
logic S_s6_291, C_s6_291;
FA FA_s6_291(.A(S_s7_295), .B(S_s7_294), .c_in(S_s7_293), .S(S_s6_291), .c_out(C_s6_291));
logic S_s6_292, C_s6_292;
FA FA_s6_292(.A(S_s7_292), .B(S_s7_291), .c_in(S_s7_290), .S(S_s6_292), .c_out(C_s6_292));
logic S_s6_293, C_s6_293;
FA FA_s6_293(.A(C_s7_288), .B(C_s7_287), .c_in(C_s7_286), .S(S_s6_293), .c_out(C_s6_293));
logic S_s6_294, C_s6_294;
FA FA_s6_294(.A(C_s7_285), .B(C_s7_284), .c_in(C_s7_283), .S(S_s6_294), .c_out(C_s6_294));
logic S_s6_295, C_s6_295;
FA FA_s6_295(.A(C_s7_282), .B(C_s7_281), .c_in(C_s7_280), .S(S_s6_295), .c_out(C_s6_295));
logic S_s6_300, C_s6_300;
FA FA_s6_300(.A(S_s7_308), .B(S_s7_307), .c_in(S_s7_306), .S(S_s6_300), .c_out(C_s6_300));
logic S_s6_301, C_s6_301;
FA FA_s6_301(.A(S_s7_305), .B(S_s7_304), .c_in(S_s7_303), .S(S_s6_301), .c_out(C_s6_301));
logic S_s6_302, C_s6_302;
FA FA_s6_302(.A(S_s7_302), .B(S_s7_301), .c_in(S_s7_300), .S(S_s6_302), .c_out(C_s6_302));
logic S_s6_303, C_s6_303;
FA FA_s6_303(.A(C_s7_298), .B(C_s7_297), .c_in(C_s7_296), .S(S_s6_303), .c_out(C_s6_303));
logic S_s6_304, C_s6_304;
FA FA_s6_304(.A(C_s7_295), .B(C_s7_294), .c_in(C_s7_293), .S(S_s6_304), .c_out(C_s6_304));
logic S_s6_305, C_s6_305;
FA FA_s6_305(.A(C_s7_292), .B(C_s7_291), .c_in(C_s7_290), .S(S_s6_305), .c_out(C_s6_305));
logic S_s6_310, C_s6_310;
FA FA_s6_310(.A(S_s7_318), .B(S_s7_317), .c_in(S_s7_316), .S(S_s6_310), .c_out(C_s6_310));
logic S_s6_311, C_s6_311;
FA FA_s6_311(.A(S_s7_315), .B(S_s7_314), .c_in(S_s7_313), .S(S_s6_311), .c_out(C_s6_311));
logic S_s6_312, C_s6_312;
FA FA_s6_312(.A(S_s7_312), .B(S_s7_311), .c_in(S_s7_310), .S(S_s6_312), .c_out(C_s6_312));
logic S_s6_313, C_s6_313;
FA FA_s6_313(.A(C_s7_308), .B(C_s7_307), .c_in(C_s7_306), .S(S_s6_313), .c_out(C_s6_313));
logic S_s6_314, C_s6_314;
FA FA_s6_314(.A(C_s7_305), .B(C_s7_304), .c_in(C_s7_303), .S(S_s6_314), .c_out(C_s6_314));
logic S_s6_315, C_s6_315;
FA FA_s6_315(.A(C_s7_302), .B(C_s7_301), .c_in(C_s7_300), .S(S_s6_315), .c_out(C_s6_315));
logic S_s6_320, C_s6_320;
FA FA_s6_320(.A(S_s7_328), .B(S_s7_327), .c_in(S_s7_326), .S(S_s6_320), .c_out(C_s6_320));
logic S_s6_321, C_s6_321;
FA FA_s6_321(.A(S_s7_325), .B(S_s7_324), .c_in(S_s7_323), .S(S_s6_321), .c_out(C_s6_321));
logic S_s6_322, C_s6_322;
FA FA_s6_322(.A(S_s7_322), .B(S_s7_321), .c_in(S_s7_320), .S(S_s6_322), .c_out(C_s6_322));
logic S_s6_323, C_s6_323;
FA FA_s6_323(.A(C_s7_318), .B(C_s7_317), .c_in(C_s7_316), .S(S_s6_323), .c_out(C_s6_323));
logic S_s6_324, C_s6_324;
FA FA_s6_324(.A(C_s7_315), .B(C_s7_314), .c_in(C_s7_313), .S(S_s6_324), .c_out(C_s6_324));
logic S_s6_325, C_s6_325;
FA FA_s6_325(.A(C_s7_312), .B(C_s7_311), .c_in(C_s7_310), .S(S_s6_325), .c_out(C_s6_325));
logic S_s6_330, C_s6_330;
FA FA_s6_330(.A(S_s7_338), .B(S_s7_337), .c_in(S_s7_336), .S(S_s6_330), .c_out(C_s6_330));
logic S_s6_331, C_s6_331;
FA FA_s6_331(.A(S_s7_335), .B(S_s7_334), .c_in(S_s7_333), .S(S_s6_331), .c_out(C_s6_331));
logic S_s6_332, C_s6_332;
FA FA_s6_332(.A(S_s7_332), .B(S_s7_331), .c_in(S_s7_330), .S(S_s6_332), .c_out(C_s6_332));
logic S_s6_333, C_s6_333;
FA FA_s6_333(.A(C_s7_328), .B(C_s7_327), .c_in(C_s7_326), .S(S_s6_333), .c_out(C_s6_333));
logic S_s6_334, C_s6_334;
FA FA_s6_334(.A(C_s7_325), .B(C_s7_324), .c_in(C_s7_323), .S(S_s6_334), .c_out(C_s6_334));
logic S_s6_335, C_s6_335;
FA FA_s6_335(.A(C_s7_322), .B(C_s7_321), .c_in(C_s7_320), .S(S_s6_335), .c_out(C_s6_335));
logic S_s6_340, C_s6_340;
FA FA_s6_340(.A(S_s7_348), .B(S_s7_347), .c_in(S_s7_346), .S(S_s6_340), .c_out(C_s6_340));
logic S_s6_341, C_s6_341;
FA FA_s6_341(.A(S_s7_345), .B(S_s7_344), .c_in(S_s7_343), .S(S_s6_341), .c_out(C_s6_341));
logic S_s6_342, C_s6_342;
FA FA_s6_342(.A(S_s7_342), .B(S_s7_341), .c_in(S_s7_340), .S(S_s6_342), .c_out(C_s6_342));
logic S_s6_343, C_s6_343;
FA FA_s6_343(.A(C_s7_338), .B(C_s7_337), .c_in(C_s7_336), .S(S_s6_343), .c_out(C_s6_343));
logic S_s6_344, C_s6_344;
FA FA_s6_344(.A(C_s7_335), .B(C_s7_334), .c_in(C_s7_333), .S(S_s6_344), .c_out(C_s6_344));
logic S_s6_345, C_s6_345;
FA FA_s6_345(.A(C_s7_332), .B(C_s7_331), .c_in(C_s7_330), .S(S_s6_345), .c_out(C_s6_345));
logic S_s6_350, C_s6_350;
FA FA_s6_350(.A(S_s7_358), .B(S_s7_357), .c_in(S_s7_356), .S(S_s6_350), .c_out(C_s6_350));
logic S_s6_351, C_s6_351;
FA FA_s6_351(.A(S_s7_355), .B(S_s7_354), .c_in(S_s7_353), .S(S_s6_351), .c_out(C_s6_351));
logic S_s6_352, C_s6_352;
FA FA_s6_352(.A(S_s7_352), .B(S_s7_351), .c_in(S_s7_350), .S(S_s6_352), .c_out(C_s6_352));
logic S_s6_353, C_s6_353;
FA FA_s6_353(.A(C_s7_348), .B(C_s7_347), .c_in(C_s7_346), .S(S_s6_353), .c_out(C_s6_353));
logic S_s6_354, C_s6_354;
FA FA_s6_354(.A(C_s7_345), .B(C_s7_344), .c_in(C_s7_343), .S(S_s6_354), .c_out(C_s6_354));
logic S_s6_355, C_s6_355;
FA FA_s6_355(.A(C_s7_342), .B(C_s7_341), .c_in(C_s7_340), .S(S_s6_355), .c_out(C_s6_355));
logic S_s6_360, C_s6_360;
FA FA_s6_360(.A(S_s7_368), .B(S_s7_367), .c_in(S_s7_366), .S(S_s6_360), .c_out(C_s6_360));
logic S_s6_361, C_s6_361;
FA FA_s6_361(.A(S_s7_365), .B(S_s7_364), .c_in(S_s7_363), .S(S_s6_361), .c_out(C_s6_361));
logic S_s6_362, C_s6_362;
FA FA_s6_362(.A(S_s7_362), .B(S_s7_361), .c_in(S_s7_360), .S(S_s6_362), .c_out(C_s6_362));
logic S_s6_363, C_s6_363;
FA FA_s6_363(.A(C_s7_358), .B(C_s7_357), .c_in(C_s7_356), .S(S_s6_363), .c_out(C_s6_363));
logic S_s6_364, C_s6_364;
FA FA_s6_364(.A(C_s7_355), .B(C_s7_354), .c_in(C_s7_353), .S(S_s6_364), .c_out(C_s6_364));
logic S_s6_365, C_s6_365;
FA FA_s6_365(.A(C_s7_352), .B(C_s7_351), .c_in(C_s7_350), .S(S_s6_365), .c_out(C_s6_365));
logic S_s6_370, C_s6_370;
FA FA_s6_370(.A(S_s7_377), .B(S_s7_376), .c_in(S_s7_375), .S(S_s6_370), .c_out(C_s6_370));
logic S_s6_371, C_s6_371;
FA FA_s6_371(.A(S_s7_374), .B(S_s7_373), .c_in(S_s7_372), .S(S_s6_371), .c_out(C_s6_371));
logic S_s6_372, C_s6_372;
FA FA_s6_372(.A(S_s7_371), .B(S_s7_370), .c_in(C_s7_368), .S(S_s6_372), .c_out(C_s6_372));
logic S_s6_373, C_s6_373;
FA FA_s6_373(.A(C_s7_367), .B(C_s7_366), .c_in(C_s7_365), .S(S_s6_373), .c_out(C_s6_373));
logic S_s6_374, C_s6_374;
FA FA_s6_374(.A(C_s7_364), .B(C_s7_363), .c_in(C_s7_362), .S(S_s6_374), .c_out(C_s6_374));
logic S_s6_375, C_s6_375;
FA FA_s6_375(.A(C_s7_361), .B(C_s7_360), .c_in(comb[30][7]), .S(S_s6_375), .c_out(C_s6_375));
logic S_s6_380, C_s6_380;
FA FA_s6_380(.A(S_s7_386), .B(S_s7_385), .c_in(S_s7_384), .S(S_s6_380), .c_out(C_s6_380));
logic S_s6_381, C_s6_381;
FA FA_s6_381(.A(S_s7_383), .B(S_s7_382), .c_in(S_s7_381), .S(S_s6_381), .c_out(C_s6_381));
logic S_s6_382, C_s6_382;
FA FA_s6_382(.A(S_s7_380), .B(C_s7_377), .c_in(C_s7_376), .S(S_s6_382), .c_out(C_s6_382));
logic S_s6_383, C_s6_383;
FA FA_s6_383(.A(C_s7_375), .B(C_s7_374), .c_in(C_s7_373), .S(S_s6_383), .c_out(C_s6_383));
logic S_s6_384, C_s6_384;
FA FA_s6_384(.A(C_s7_372), .B(C_s7_371), .c_in(C_s7_370), .S(S_s6_384), .c_out(C_s6_384));
logic S_s6_385, C_s6_385;
FA FA_s6_385(.A(comb[28][10]), .B(comb[29][9]), .c_in(comb[30][8]), .S(S_s6_385), .c_out(C_s6_385));
logic S_s6_390, C_s6_390;
FA FA_s6_390(.A(S_s7_395), .B(S_s7_394), .c_in(S_s7_393), .S(S_s6_390), .c_out(C_s6_390));
logic S_s6_391, C_s6_391;
FA FA_s6_391(.A(S_s7_392), .B(S_s7_391), .c_in(S_s7_390), .S(S_s6_391), .c_out(C_s6_391));
logic S_s6_392, C_s6_392;
FA FA_s6_392(.A(C_s7_386), .B(C_s7_385), .c_in(C_s7_384), .S(S_s6_392), .c_out(C_s6_392));
logic S_s6_393, C_s6_393;
FA FA_s6_393(.A(C_s7_383), .B(C_s7_382), .c_in(C_s7_381), .S(S_s6_393), .c_out(C_s6_393));
logic S_s6_394, C_s6_394;
FA FA_s6_394(.A(C_s7_380), .B(comb[26][13]), .c_in(comb[27][12]), .S(S_s6_394), .c_out(C_s6_394));
logic S_s6_395, C_s6_395;
FA FA_s6_395(.A(comb[28][11]), .B(comb[29][10]), .c_in(comb[30][9]), .S(S_s6_395), .c_out(C_s6_395));
logic S_s6_400, C_s6_400;
FA FA_s6_400(.A(S_s7_404), .B(S_s7_403), .c_in(S_s7_402), .S(S_s6_400), .c_out(C_s6_400));
logic S_s6_401, C_s6_401;
FA FA_s6_401(.A(S_s7_401), .B(S_s7_400), .c_in(C_s7_395), .S(S_s6_401), .c_out(C_s6_401));
logic S_s6_402, C_s6_402;
FA FA_s6_402(.A(C_s7_394), .B(C_s7_393), .c_in(C_s7_392), .S(S_s6_402), .c_out(C_s6_402));
logic S_s6_403, C_s6_403;
FA FA_s6_403(.A(C_s7_391), .B(C_s7_390), .c_in(comb[24][16]), .S(S_s6_403), .c_out(C_s6_403));
logic S_s6_404, C_s6_404;
FA FA_s6_404(.A(comb[25][15]), .B(comb[26][14]), .c_in(comb[27][13]), .S(S_s6_404), .c_out(C_s6_404));
logic S_s6_405, C_s6_405;
FA FA_s6_405(.A(comb[28][12]), .B(comb[29][11]), .c_in(comb[30][10]), .S(S_s6_405), .c_out(C_s6_405));
logic S_s6_410, C_s6_410;
FA FA_s6_410(.A(S_s7_413), .B(S_s7_412), .c_in(S_s7_411), .S(S_s6_410), .c_out(C_s6_410));
logic S_s6_411, C_s6_411;
FA FA_s6_411(.A(S_s7_410), .B(C_s7_404), .c_in(C_s7_403), .S(S_s6_411), .c_out(C_s6_411));
logic S_s6_412, C_s6_412;
FA FA_s6_412(.A(C_s7_402), .B(C_s7_401), .c_in(C_s7_400), .S(S_s6_412), .c_out(C_s6_412));
logic S_s6_413, C_s6_413;
FA FA_s6_413(.A(comb[22][19]), .B(comb[23][18]), .c_in(comb[24][17]), .S(S_s6_413), .c_out(C_s6_413));
logic S_s6_414, C_s6_414;
FA FA_s6_414(.A(comb[25][16]), .B(comb[26][15]), .c_in(comb[27][14]), .S(S_s6_414), .c_out(C_s6_414));
logic S_s6_415, C_s6_415;
FA FA_s6_415(.A(comb[28][13]), .B(comb[29][12]), .c_in(comb[30][11]), .S(S_s6_415), .c_out(C_s6_415));
logic S_s6_420, C_s6_420;
FA FA_s6_420(.A(S_s7_422), .B(S_s7_421), .c_in(S_s7_420), .S(S_s6_420), .c_out(C_s6_420));
logic S_s6_421, C_s6_421;
FA FA_s6_421(.A(C_s7_413), .B(C_s7_412), .c_in(C_s7_411), .S(S_s6_421), .c_out(C_s6_421));
logic S_s6_422, C_s6_422;
FA FA_s6_422(.A(C_s7_410), .B(comb[20][22]), .c_in(comb[21][21]), .S(S_s6_422), .c_out(C_s6_422));
logic S_s6_423, C_s6_423;
FA FA_s6_423(.A(comb[22][20]), .B(comb[23][19]), .c_in(comb[24][18]), .S(S_s6_423), .c_out(C_s6_423));
logic S_s6_424, C_s6_424;
FA FA_s6_424(.A(comb[25][17]), .B(comb[26][16]), .c_in(comb[27][15]), .S(S_s6_424), .c_out(C_s6_424));
logic S_s6_425, C_s6_425;
FA FA_s6_425(.A(comb[28][14]), .B(comb[29][13]), .c_in(comb[30][12]), .S(S_s6_425), .c_out(C_s6_425));
logic S_s6_430, C_s6_430;
FA FA_s6_430(.A(S_s7_431), .B(S_s7_430), .c_in(C_s7_422), .S(S_s6_430), .c_out(C_s6_430));
logic S_s6_431, C_s6_431;
FA FA_s6_431(.A(C_s7_421), .B(C_s7_420), .c_in(comb[18][25]), .S(S_s6_431), .c_out(C_s6_431));
logic S_s6_432, C_s6_432;
FA FA_s6_432(.A(comb[19][24]), .B(comb[20][23]), .c_in(comb[21][22]), .S(S_s6_432), .c_out(C_s6_432));
logic S_s6_433, C_s6_433;
FA FA_s6_433(.A(comb[22][21]), .B(comb[23][20]), .c_in(comb[24][19]), .S(S_s6_433), .c_out(C_s6_433));
logic S_s6_434, C_s6_434;
FA FA_s6_434(.A(comb[25][18]), .B(comb[26][17]), .c_in(comb[27][16]), .S(S_s6_434), .c_out(C_s6_434));
logic S_s6_435, C_s6_435;
FA FA_s6_435(.A(comb[28][15]), .B(comb[29][14]), .c_in(comb[30][13]), .S(S_s6_435), .c_out(C_s6_435));
logic S_s6_440, C_s6_440;
FA FA_s6_440(.A(S_s7_440), .B(C_s7_431), .c_in(C_s7_430), .S(S_s6_440), .c_out(C_s6_440));
logic S_s6_441, C_s6_441;
FA FA_s6_441(.A(comb[16][28]), .B(comb[17][27]), .c_in(comb[18][26]), .S(S_s6_441), .c_out(C_s6_441));
logic S_s6_442, C_s6_442;
FA FA_s6_442(.A(comb[19][25]), .B(comb[20][24]), .c_in(comb[21][23]), .S(S_s6_442), .c_out(C_s6_442));
logic S_s6_443, C_s6_443;
FA FA_s6_443(.A(comb[22][22]), .B(comb[23][21]), .c_in(comb[24][20]), .S(S_s6_443), .c_out(C_s6_443));
logic S_s6_444, C_s6_444;
FA FA_s6_444(.A(comb[25][19]), .B(comb[26][18]), .c_in(comb[27][17]), .S(S_s6_444), .c_out(C_s6_444));
logic S_s6_445, C_s6_445;
FA FA_s6_445(.A(comb[28][16]), .B(comb[29][15]), .c_in(comb[30][14]), .S(S_s6_445), .c_out(C_s6_445));
logic S_s6_450, C_s6_450;
FA FA_s6_450(.A(C_s7_440), .B(comb[14][31]), .c_in(comb[15][30]), .S(S_s6_450), .c_out(C_s6_450));
logic S_s6_451, C_s6_451;
FA FA_s6_451(.A(comb[16][29]), .B(comb[17][28]), .c_in(comb[18][27]), .S(S_s6_451), .c_out(C_s6_451));
logic S_s6_452, C_s6_452;
FA FA_s6_452(.A(comb[19][26]), .B(comb[20][25]), .c_in(comb[21][24]), .S(S_s6_452), .c_out(C_s6_452));
logic S_s6_453, C_s6_453;
FA FA_s6_453(.A(comb[22][23]), .B(comb[23][22]), .c_in(comb[24][21]), .S(S_s6_453), .c_out(C_s6_453));
logic S_s6_454, C_s6_454;
FA FA_s6_454(.A(comb[25][20]), .B(comb[26][19]), .c_in(comb[27][18]), .S(S_s6_454), .c_out(C_s6_454));
logic S_s6_455, C_s6_455;
FA FA_s6_455(.A(comb[28][17]), .B(comb[29][16]), .c_in(comb[30][15]), .S(S_s6_455), .c_out(C_s6_455));
logic S_s6_460, C_s6_460;
FA FA_s6_460(.A(comb[15][31]), .B(comb[16][30]), .c_in(comb[17][29]), .S(S_s6_460), .c_out(C_s6_460));
logic S_s6_461, C_s6_461;
FA FA_s6_461(.A(comb[18][28]), .B(comb[19][27]), .c_in(comb[20][26]), .S(S_s6_461), .c_out(C_s6_461));
logic S_s6_462, C_s6_462;
FA FA_s6_462(.A(comb[21][25]), .B(comb[22][24]), .c_in(comb[23][23]), .S(S_s6_462), .c_out(C_s6_462));
logic S_s6_463, C_s6_463;
FA FA_s6_463(.A(comb[24][22]), .B(comb[25][21]), .c_in(comb[26][20]), .S(S_s6_463), .c_out(C_s6_463));
logic S_s6_464, C_s6_464;
FA FA_s6_464(.A(comb[27][19]), .B(comb[28][18]), .c_in(comb[29][17]), .S(S_s6_464), .c_out(C_s6_464));
logic S_s6_470, C_s6_470;
FA FA_s6_470(.A(comb[16][31]), .B(comb[17][30]), .c_in(comb[18][29]), .S(S_s6_470), .c_out(C_s6_470));
logic S_s6_471, C_s6_471;
FA FA_s6_471(.A(comb[19][28]), .B(comb[20][27]), .c_in(comb[21][26]), .S(S_s6_471), .c_out(C_s6_471));
logic S_s6_472, C_s6_472;
FA FA_s6_472(.A(comb[22][25]), .B(comb[23][24]), .c_in(comb[24][23]), .S(S_s6_472), .c_out(C_s6_472));
logic S_s6_473, C_s6_473;
FA FA_s6_473(.A(comb[25][22]), .B(comb[26][21]), .c_in(comb[27][20]), .S(S_s6_473), .c_out(C_s6_473));
logic S_s6_480, C_s6_480;
FA FA_s6_480(.A(comb[17][31]), .B(comb[18][30]), .c_in(comb[19][29]), .S(S_s6_480), .c_out(C_s6_480));
logic S_s6_481, C_s6_481;
FA FA_s6_481(.A(comb[20][28]), .B(comb[21][27]), .c_in(comb[22][26]), .S(S_s6_481), .c_out(C_s6_481));
logic S_s6_482, C_s6_482;
FA FA_s6_482(.A(comb[23][25]), .B(comb[24][24]), .c_in(comb[25][23]), .S(S_s6_482), .c_out(C_s6_482));
logic S_s6_490, C_s6_490;
FA FA_s6_490(.A(comb[18][31]), .B(comb[19][30]), .c_in(comb[20][29]), .S(S_s6_490), .c_out(C_s6_490));
logic S_s6_491, C_s6_491;
FA FA_s6_491(.A(comb[21][28]), .B(comb[22][27]), .c_in(comb[23][26]), .S(S_s6_491), .c_out(C_s6_491));
logic S_s6_500, C_s6_500;
FA FA_s6_500(.A(comb[19][31]), .B(comb[20][30]), .c_in(comb[21][29]), .S(S_s6_500), .c_out(C_s6_500));
// stage 6 end ======================================================================================================= 

// stage 5 begin ======================================================================================================= 
logic S_s5_90, C_s5_90;
HA HA_s5_90(.A(comb[0][9]), .B(comb[1][8]), .S(S_s5_90), .c_out(C_s5_90));
logic S_s5_100, C_s5_100;
FA FA_s5_100(.A(comb[0][10]), .B(comb[1][9]), .c_in(comb[2][8]), .S(S_s5_100), .c_out(C_s5_100));
logic S_s5_101, C_s5_101;
HA HA_s5_101(.A(comb[3][7]), .B(comb[4][6]), .S(S_s5_101), .c_out(C_s5_101));
logic S_s5_110, C_s5_110;
FA FA_s5_110(.A(comb[0][11]), .B(comb[1][10]), .c_in(comb[2][9]), .S(S_s5_110), .c_out(C_s5_110));
logic S_s5_111, C_s5_111;
FA FA_s5_111(.A(comb[3][8]), .B(comb[4][7]), .c_in(comb[5][6]), .S(S_s5_111), .c_out(C_s5_111));
logic S_s5_112, C_s5_112;
HA HA_s5_112(.A(comb[6][5]), .B(comb[7][4]), .S(S_s5_112), .c_out(C_s5_112));
logic S_s5_120, C_s5_120;
FA FA_s5_120(.A(comb[0][12]), .B(comb[1][11]), .c_in(comb[2][10]), .S(S_s5_120), .c_out(C_s5_120));
logic S_s5_121, C_s5_121;
FA FA_s5_121(.A(comb[3][9]), .B(comb[4][8]), .c_in(comb[5][7]), .S(S_s5_121), .c_out(C_s5_121));
logic S_s5_122, C_s5_122;
FA FA_s5_122(.A(comb[6][6]), .B(comb[7][5]), .c_in(comb[8][4]), .S(S_s5_122), .c_out(C_s5_122));
logic S_s5_123, C_s5_123;
HA HA_s5_123(.A(comb[9][3]), .B(comb[10][2]), .S(S_s5_123), .c_out(C_s5_123));
logic S_s5_130, C_s5_130;
FA FA_s5_130(.A(S_s6_130), .B(comb[2][11]), .c_in(comb[3][10]), .S(S_s5_130), .c_out(C_s5_130));
logic S_s5_131, C_s5_131;
FA FA_s5_131(.A(comb[4][9]), .B(comb[5][8]), .c_in(comb[6][7]), .S(S_s5_131), .c_out(C_s5_131));
logic S_s5_132, C_s5_132;
FA FA_s5_132(.A(comb[7][6]), .B(comb[8][5]), .c_in(comb[9][4]), .S(S_s5_132), .c_out(C_s5_132));
logic S_s5_133, C_s5_133;
FA FA_s5_133(.A(comb[10][3]), .B(comb[11][2]), .c_in(comb[12][1]), .S(S_s5_133), .c_out(C_s5_133));
logic S_s5_140, C_s5_140;
FA FA_s5_140(.A(S_s6_141), .B(S_s6_140), .c_in(C_s6_130), .S(S_s5_140), .c_out(C_s5_140));
logic S_s5_141, C_s5_141;
FA FA_s5_141(.A(comb[5][9]), .B(comb[6][8]), .c_in(comb[7][7]), .S(S_s5_141), .c_out(C_s5_141));
logic S_s5_142, C_s5_142;
FA FA_s5_142(.A(comb[8][6]), .B(comb[9][5]), .c_in(comb[10][4]), .S(S_s5_142), .c_out(C_s5_142));
logic S_s5_143, C_s5_143;
FA FA_s5_143(.A(comb[11][3]), .B(comb[12][2]), .c_in(comb[13][1]), .S(S_s5_143), .c_out(C_s5_143));
logic S_s5_150, C_s5_150;
FA FA_s5_150(.A(S_s6_152), .B(S_s6_151), .c_in(S_s6_150), .S(S_s5_150), .c_out(C_s5_150));
logic S_s5_151, C_s5_151;
FA FA_s5_151(.A(C_s6_141), .B(C_s6_140), .c_in(comb[8][7]), .S(S_s5_151), .c_out(C_s5_151));
logic S_s5_152, C_s5_152;
FA FA_s5_152(.A(comb[9][6]), .B(comb[10][5]), .c_in(comb[11][4]), .S(S_s5_152), .c_out(C_s5_152));
logic S_s5_153, C_s5_153;
FA FA_s5_153(.A(comb[12][3]), .B(comb[13][2]), .c_in(comb[14][1]), .S(S_s5_153), .c_out(C_s5_153));
logic S_s5_160, C_s5_160;
FA FA_s5_160(.A(S_s6_163), .B(S_s6_162), .c_in(S_s6_161), .S(S_s5_160), .c_out(C_s5_160));
logic S_s5_161, C_s5_161;
FA FA_s5_161(.A(S_s6_160), .B(C_s6_152), .c_in(C_s6_151), .S(S_s5_161), .c_out(C_s5_161));
logic S_s5_162, C_s5_162;
FA FA_s5_162(.A(C_s6_150), .B(comb[11][5]), .c_in(comb[12][4]), .S(S_s5_162), .c_out(C_s5_162));
logic S_s5_163, C_s5_163;
FA FA_s5_163(.A(comb[13][3]), .B(comb[14][2]), .c_in(comb[15][1]), .S(S_s5_163), .c_out(C_s5_163));
logic S_s5_170, C_s5_170;
FA FA_s5_170(.A(S_s6_174), .B(S_s6_173), .c_in(S_s6_172), .S(S_s5_170), .c_out(C_s5_170));
logic S_s5_171, C_s5_171;
FA FA_s5_171(.A(S_s6_171), .B(S_s6_170), .c_in(C_s6_163), .S(S_s5_171), .c_out(C_s5_171));
logic S_s5_172, C_s5_172;
FA FA_s5_172(.A(C_s6_162), .B(C_s6_161), .c_in(C_s6_160), .S(S_s5_172), .c_out(C_s5_172));
logic S_s5_173, C_s5_173;
FA FA_s5_173(.A(comb[14][3]), .B(comb[15][2]), .c_in(comb[16][1]), .S(S_s5_173), .c_out(C_s5_173));
logic S_s5_180, C_s5_180;
FA FA_s5_180(.A(S_s6_185), .B(S_s6_184), .c_in(S_s6_183), .S(S_s5_180), .c_out(C_s5_180));
logic S_s5_181, C_s5_181;
FA FA_s5_181(.A(S_s6_182), .B(S_s6_181), .c_in(S_s6_180), .S(S_s5_181), .c_out(C_s5_181));
logic S_s5_182, C_s5_182;
FA FA_s5_182(.A(C_s6_174), .B(C_s6_173), .c_in(C_s6_172), .S(S_s5_182), .c_out(C_s5_182));
logic S_s5_183, C_s5_183;
FA FA_s5_183(.A(C_s6_171), .B(C_s6_170), .c_in(comb[17][1]), .S(S_s5_183), .c_out(C_s5_183));
logic S_s5_190, C_s5_190;
FA FA_s5_190(.A(S_s6_195), .B(S_s6_194), .c_in(S_s6_193), .S(S_s5_190), .c_out(C_s5_190));
logic S_s5_191, C_s5_191;
FA FA_s5_191(.A(S_s6_192), .B(S_s6_191), .c_in(S_s6_190), .S(S_s5_191), .c_out(C_s5_191));
logic S_s5_192, C_s5_192;
FA FA_s5_192(.A(C_s6_185), .B(C_s6_184), .c_in(C_s6_183), .S(S_s5_192), .c_out(C_s5_192));
logic S_s5_193, C_s5_193;
FA FA_s5_193(.A(C_s6_182), .B(C_s6_181), .c_in(C_s6_180), .S(S_s5_193), .c_out(C_s5_193));
logic S_s5_200, C_s5_200;
FA FA_s5_200(.A(S_s6_205), .B(S_s6_204), .c_in(S_s6_203), .S(S_s5_200), .c_out(C_s5_200));
logic S_s5_201, C_s5_201;
FA FA_s5_201(.A(S_s6_202), .B(S_s6_201), .c_in(S_s6_200), .S(S_s5_201), .c_out(C_s5_201));
logic S_s5_202, C_s5_202;
FA FA_s5_202(.A(C_s6_195), .B(C_s6_194), .c_in(C_s6_193), .S(S_s5_202), .c_out(C_s5_202));
logic S_s5_203, C_s5_203;
FA FA_s5_203(.A(C_s6_192), .B(C_s6_191), .c_in(C_s6_190), .S(S_s5_203), .c_out(C_s5_203));
logic S_s5_210, C_s5_210;
FA FA_s5_210(.A(S_s6_215), .B(S_s6_214), .c_in(S_s6_213), .S(S_s5_210), .c_out(C_s5_210));
logic S_s5_211, C_s5_211;
FA FA_s5_211(.A(S_s6_212), .B(S_s6_211), .c_in(S_s6_210), .S(S_s5_211), .c_out(C_s5_211));
logic S_s5_212, C_s5_212;
FA FA_s5_212(.A(C_s6_205), .B(C_s6_204), .c_in(C_s6_203), .S(S_s5_212), .c_out(C_s5_212));
logic S_s5_213, C_s5_213;
FA FA_s5_213(.A(C_s6_202), .B(C_s6_201), .c_in(C_s6_200), .S(S_s5_213), .c_out(C_s5_213));
logic S_s5_220, C_s5_220;
FA FA_s5_220(.A(S_s6_225), .B(S_s6_224), .c_in(S_s6_223), .S(S_s5_220), .c_out(C_s5_220));
logic S_s5_221, C_s5_221;
FA FA_s5_221(.A(S_s6_222), .B(S_s6_221), .c_in(S_s6_220), .S(S_s5_221), .c_out(C_s5_221));
logic S_s5_222, C_s5_222;
FA FA_s5_222(.A(C_s6_215), .B(C_s6_214), .c_in(C_s6_213), .S(S_s5_222), .c_out(C_s5_222));
logic S_s5_223, C_s5_223;
FA FA_s5_223(.A(C_s6_212), .B(C_s6_211), .c_in(C_s6_210), .S(S_s5_223), .c_out(C_s5_223));
logic S_s5_230, C_s5_230;
FA FA_s5_230(.A(S_s6_235), .B(S_s6_234), .c_in(S_s6_233), .S(S_s5_230), .c_out(C_s5_230));
logic S_s5_231, C_s5_231;
FA FA_s5_231(.A(S_s6_232), .B(S_s6_231), .c_in(S_s6_230), .S(S_s5_231), .c_out(C_s5_231));
logic S_s5_232, C_s5_232;
FA FA_s5_232(.A(C_s6_225), .B(C_s6_224), .c_in(C_s6_223), .S(S_s5_232), .c_out(C_s5_232));
logic S_s5_233, C_s5_233;
FA FA_s5_233(.A(C_s6_222), .B(C_s6_221), .c_in(C_s6_220), .S(S_s5_233), .c_out(C_s5_233));
logic S_s5_240, C_s5_240;
FA FA_s5_240(.A(S_s6_245), .B(S_s6_244), .c_in(S_s6_243), .S(S_s5_240), .c_out(C_s5_240));
logic S_s5_241, C_s5_241;
FA FA_s5_241(.A(S_s6_242), .B(S_s6_241), .c_in(S_s6_240), .S(S_s5_241), .c_out(C_s5_241));
logic S_s5_242, C_s5_242;
FA FA_s5_242(.A(C_s6_235), .B(C_s6_234), .c_in(C_s6_233), .S(S_s5_242), .c_out(C_s5_242));
logic S_s5_243, C_s5_243;
FA FA_s5_243(.A(C_s6_232), .B(C_s6_231), .c_in(C_s6_230), .S(S_s5_243), .c_out(C_s5_243));
logic S_s5_250, C_s5_250;
FA FA_s5_250(.A(S_s6_255), .B(S_s6_254), .c_in(S_s6_253), .S(S_s5_250), .c_out(C_s5_250));
logic S_s5_251, C_s5_251;
FA FA_s5_251(.A(S_s6_252), .B(S_s6_251), .c_in(S_s6_250), .S(S_s5_251), .c_out(C_s5_251));
logic S_s5_252, C_s5_252;
FA FA_s5_252(.A(C_s6_245), .B(C_s6_244), .c_in(C_s6_243), .S(S_s5_252), .c_out(C_s5_252));
logic S_s5_253, C_s5_253;
FA FA_s5_253(.A(C_s6_242), .B(C_s6_241), .c_in(C_s6_240), .S(S_s5_253), .c_out(C_s5_253));
logic S_s5_260, C_s5_260;
FA FA_s5_260(.A(S_s6_265), .B(S_s6_264), .c_in(S_s6_263), .S(S_s5_260), .c_out(C_s5_260));
logic S_s5_261, C_s5_261;
FA FA_s5_261(.A(S_s6_262), .B(S_s6_261), .c_in(S_s6_260), .S(S_s5_261), .c_out(C_s5_261));
logic S_s5_262, C_s5_262;
FA FA_s5_262(.A(C_s6_255), .B(C_s6_254), .c_in(C_s6_253), .S(S_s5_262), .c_out(C_s5_262));
logic S_s5_263, C_s5_263;
FA FA_s5_263(.A(C_s6_252), .B(C_s6_251), .c_in(C_s6_250), .S(S_s5_263), .c_out(C_s5_263));
logic S_s5_270, C_s5_270;
FA FA_s5_270(.A(S_s6_275), .B(S_s6_274), .c_in(S_s6_273), .S(S_s5_270), .c_out(C_s5_270));
logic S_s5_271, C_s5_271;
FA FA_s5_271(.A(S_s6_272), .B(S_s6_271), .c_in(S_s6_270), .S(S_s5_271), .c_out(C_s5_271));
logic S_s5_272, C_s5_272;
FA FA_s5_272(.A(C_s6_265), .B(C_s6_264), .c_in(C_s6_263), .S(S_s5_272), .c_out(C_s5_272));
logic S_s5_273, C_s5_273;
FA FA_s5_273(.A(C_s6_262), .B(C_s6_261), .c_in(C_s6_260), .S(S_s5_273), .c_out(C_s5_273));
logic S_s5_280, C_s5_280;
FA FA_s5_280(.A(S_s6_285), .B(S_s6_284), .c_in(S_s6_283), .S(S_s5_280), .c_out(C_s5_280));
logic S_s5_281, C_s5_281;
FA FA_s5_281(.A(S_s6_282), .B(S_s6_281), .c_in(S_s6_280), .S(S_s5_281), .c_out(C_s5_281));
logic S_s5_282, C_s5_282;
FA FA_s5_282(.A(C_s6_275), .B(C_s6_274), .c_in(C_s6_273), .S(S_s5_282), .c_out(C_s5_282));
logic S_s5_283, C_s5_283;
FA FA_s5_283(.A(C_s6_272), .B(C_s6_271), .c_in(C_s6_270), .S(S_s5_283), .c_out(C_s5_283));
logic S_s5_290, C_s5_290;
FA FA_s5_290(.A(S_s6_295), .B(S_s6_294), .c_in(S_s6_293), .S(S_s5_290), .c_out(C_s5_290));
logic S_s5_291, C_s5_291;
FA FA_s5_291(.A(S_s6_292), .B(S_s6_291), .c_in(S_s6_290), .S(S_s5_291), .c_out(C_s5_291));
logic S_s5_292, C_s5_292;
FA FA_s5_292(.A(C_s6_285), .B(C_s6_284), .c_in(C_s6_283), .S(S_s5_292), .c_out(C_s5_292));
logic S_s5_293, C_s5_293;
FA FA_s5_293(.A(C_s6_282), .B(C_s6_281), .c_in(C_s6_280), .S(S_s5_293), .c_out(C_s5_293));
logic S_s5_300, C_s5_300;
FA FA_s5_300(.A(S_s6_305), .B(S_s6_304), .c_in(S_s6_303), .S(S_s5_300), .c_out(C_s5_300));
logic S_s5_301, C_s5_301;
FA FA_s5_301(.A(S_s6_302), .B(S_s6_301), .c_in(S_s6_300), .S(S_s5_301), .c_out(C_s5_301));
logic S_s5_302, C_s5_302;
FA FA_s5_302(.A(C_s6_295), .B(C_s6_294), .c_in(C_s6_293), .S(S_s5_302), .c_out(C_s5_302));
logic S_s5_303, C_s5_303;
FA FA_s5_303(.A(C_s6_292), .B(C_s6_291), .c_in(C_s6_290), .S(S_s5_303), .c_out(C_s5_303));
logic S_s5_310, C_s5_310;
FA FA_s5_310(.A(S_s6_315), .B(S_s6_314), .c_in(S_s6_313), .S(S_s5_310), .c_out(C_s5_310));
logic S_s5_311, C_s5_311;
FA FA_s5_311(.A(S_s6_312), .B(S_s6_311), .c_in(S_s6_310), .S(S_s5_311), .c_out(C_s5_311));
logic S_s5_312, C_s5_312;
FA FA_s5_312(.A(C_s6_305), .B(C_s6_304), .c_in(C_s6_303), .S(S_s5_312), .c_out(C_s5_312));
logic S_s5_313, C_s5_313;
FA FA_s5_313(.A(C_s6_302), .B(C_s6_301), .c_in(C_s6_300), .S(S_s5_313), .c_out(C_s5_313));
logic S_s5_320, C_s5_320;
FA FA_s5_320(.A(S_s6_325), .B(S_s6_324), .c_in(S_s6_323), .S(S_s5_320), .c_out(C_s5_320));
logic S_s5_321, C_s5_321;
FA FA_s5_321(.A(S_s6_322), .B(S_s6_321), .c_in(S_s6_320), .S(S_s5_321), .c_out(C_s5_321));
logic S_s5_322, C_s5_322;
FA FA_s5_322(.A(C_s6_315), .B(C_s6_314), .c_in(C_s6_313), .S(S_s5_322), .c_out(C_s5_322));
logic S_s5_323, C_s5_323;
FA FA_s5_323(.A(C_s6_312), .B(C_s6_311), .c_in(C_s6_310), .S(S_s5_323), .c_out(C_s5_323));
logic S_s5_330, C_s5_330;
FA FA_s5_330(.A(S_s6_335), .B(S_s6_334), .c_in(S_s6_333), .S(S_s5_330), .c_out(C_s5_330));
logic S_s5_331, C_s5_331;
FA FA_s5_331(.A(S_s6_332), .B(S_s6_331), .c_in(S_s6_330), .S(S_s5_331), .c_out(C_s5_331));
logic S_s5_332, C_s5_332;
FA FA_s5_332(.A(C_s6_325), .B(C_s6_324), .c_in(C_s6_323), .S(S_s5_332), .c_out(C_s5_332));
logic S_s5_333, C_s5_333;
FA FA_s5_333(.A(C_s6_322), .B(C_s6_321), .c_in(C_s6_320), .S(S_s5_333), .c_out(C_s5_333));
logic S_s5_340, C_s5_340;
FA FA_s5_340(.A(S_s6_345), .B(S_s6_344), .c_in(S_s6_343), .S(S_s5_340), .c_out(C_s5_340));
logic S_s5_341, C_s5_341;
FA FA_s5_341(.A(S_s6_342), .B(S_s6_341), .c_in(S_s6_340), .S(S_s5_341), .c_out(C_s5_341));
logic S_s5_342, C_s5_342;
FA FA_s5_342(.A(C_s6_335), .B(C_s6_334), .c_in(C_s6_333), .S(S_s5_342), .c_out(C_s5_342));
logic S_s5_343, C_s5_343;
FA FA_s5_343(.A(C_s6_332), .B(C_s6_331), .c_in(C_s6_330), .S(S_s5_343), .c_out(C_s5_343));
logic S_s5_350, C_s5_350;
FA FA_s5_350(.A(S_s6_355), .B(S_s6_354), .c_in(S_s6_353), .S(S_s5_350), .c_out(C_s5_350));
logic S_s5_351, C_s5_351;
FA FA_s5_351(.A(S_s6_352), .B(S_s6_351), .c_in(S_s6_350), .S(S_s5_351), .c_out(C_s5_351));
logic S_s5_352, C_s5_352;
FA FA_s5_352(.A(C_s6_345), .B(C_s6_344), .c_in(C_s6_343), .S(S_s5_352), .c_out(C_s5_352));
logic S_s5_353, C_s5_353;
FA FA_s5_353(.A(C_s6_342), .B(C_s6_341), .c_in(C_s6_340), .S(S_s5_353), .c_out(C_s5_353));
logic S_s5_360, C_s5_360;
FA FA_s5_360(.A(S_s6_365), .B(S_s6_364), .c_in(S_s6_363), .S(S_s5_360), .c_out(C_s5_360));
logic S_s5_361, C_s5_361;
FA FA_s5_361(.A(S_s6_362), .B(S_s6_361), .c_in(S_s6_360), .S(S_s5_361), .c_out(C_s5_361));
logic S_s5_362, C_s5_362;
FA FA_s5_362(.A(C_s6_355), .B(C_s6_354), .c_in(C_s6_353), .S(S_s5_362), .c_out(C_s5_362));
logic S_s5_363, C_s5_363;
FA FA_s5_363(.A(C_s6_352), .B(C_s6_351), .c_in(C_s6_350), .S(S_s5_363), .c_out(C_s5_363));
logic S_s5_370, C_s5_370;
FA FA_s5_370(.A(S_s6_375), .B(S_s6_374), .c_in(S_s6_373), .S(S_s5_370), .c_out(C_s5_370));
logic S_s5_371, C_s5_371;
FA FA_s5_371(.A(S_s6_372), .B(S_s6_371), .c_in(S_s6_370), .S(S_s5_371), .c_out(C_s5_371));
logic S_s5_372, C_s5_372;
FA FA_s5_372(.A(C_s6_365), .B(C_s6_364), .c_in(C_s6_363), .S(S_s5_372), .c_out(C_s5_372));
logic S_s5_373, C_s5_373;
FA FA_s5_373(.A(C_s6_362), .B(C_s6_361), .c_in(C_s6_360), .S(S_s5_373), .c_out(C_s5_373));
logic S_s5_380, C_s5_380;
FA FA_s5_380(.A(S_s6_385), .B(S_s6_384), .c_in(S_s6_383), .S(S_s5_380), .c_out(C_s5_380));
logic S_s5_381, C_s5_381;
FA FA_s5_381(.A(S_s6_382), .B(S_s6_381), .c_in(S_s6_380), .S(S_s5_381), .c_out(C_s5_381));
logic S_s5_382, C_s5_382;
FA FA_s5_382(.A(C_s6_375), .B(C_s6_374), .c_in(C_s6_373), .S(S_s5_382), .c_out(C_s5_382));
logic S_s5_383, C_s5_383;
FA FA_s5_383(.A(C_s6_372), .B(C_s6_371), .c_in(C_s6_370), .S(S_s5_383), .c_out(C_s5_383));
logic S_s5_390, C_s5_390;
FA FA_s5_390(.A(S_s6_395), .B(S_s6_394), .c_in(S_s6_393), .S(S_s5_390), .c_out(C_s5_390));
logic S_s5_391, C_s5_391;
FA FA_s5_391(.A(S_s6_392), .B(S_s6_391), .c_in(S_s6_390), .S(S_s5_391), .c_out(C_s5_391));
logic S_s5_392, C_s5_392;
FA FA_s5_392(.A(C_s6_385), .B(C_s6_384), .c_in(C_s6_383), .S(S_s5_392), .c_out(C_s5_392));
logic S_s5_393, C_s5_393;
FA FA_s5_393(.A(C_s6_382), .B(C_s6_381), .c_in(C_s6_380), .S(S_s5_393), .c_out(C_s5_393));
logic S_s5_400, C_s5_400;
FA FA_s5_400(.A(S_s6_405), .B(S_s6_404), .c_in(S_s6_403), .S(S_s5_400), .c_out(C_s5_400));
logic S_s5_401, C_s5_401;
FA FA_s5_401(.A(S_s6_402), .B(S_s6_401), .c_in(S_s6_400), .S(S_s5_401), .c_out(C_s5_401));
logic S_s5_402, C_s5_402;
FA FA_s5_402(.A(C_s6_395), .B(C_s6_394), .c_in(C_s6_393), .S(S_s5_402), .c_out(C_s5_402));
logic S_s5_403, C_s5_403;
FA FA_s5_403(.A(C_s6_392), .B(C_s6_391), .c_in(C_s6_390), .S(S_s5_403), .c_out(C_s5_403));
logic S_s5_410, C_s5_410;
FA FA_s5_410(.A(S_s6_415), .B(S_s6_414), .c_in(S_s6_413), .S(S_s5_410), .c_out(C_s5_410));
logic S_s5_411, C_s5_411;
FA FA_s5_411(.A(S_s6_412), .B(S_s6_411), .c_in(S_s6_410), .S(S_s5_411), .c_out(C_s5_411));
logic S_s5_412, C_s5_412;
FA FA_s5_412(.A(C_s6_405), .B(C_s6_404), .c_in(C_s6_403), .S(S_s5_412), .c_out(C_s5_412));
logic S_s5_413, C_s5_413;
FA FA_s5_413(.A(C_s6_402), .B(C_s6_401), .c_in(C_s6_400), .S(S_s5_413), .c_out(C_s5_413));
logic S_s5_420, C_s5_420;
FA FA_s5_420(.A(S_s6_425), .B(S_s6_424), .c_in(S_s6_423), .S(S_s5_420), .c_out(C_s5_420));
logic S_s5_421, C_s5_421;
FA FA_s5_421(.A(S_s6_422), .B(S_s6_421), .c_in(S_s6_420), .S(S_s5_421), .c_out(C_s5_421));
logic S_s5_422, C_s5_422;
FA FA_s5_422(.A(C_s6_415), .B(C_s6_414), .c_in(C_s6_413), .S(S_s5_422), .c_out(C_s5_422));
logic S_s5_423, C_s5_423;
FA FA_s5_423(.A(C_s6_412), .B(C_s6_411), .c_in(C_s6_410), .S(S_s5_423), .c_out(C_s5_423));
logic S_s5_430, C_s5_430;
FA FA_s5_430(.A(S_s6_435), .B(S_s6_434), .c_in(S_s6_433), .S(S_s5_430), .c_out(C_s5_430));
logic S_s5_431, C_s5_431;
FA FA_s5_431(.A(S_s6_432), .B(S_s6_431), .c_in(S_s6_430), .S(S_s5_431), .c_out(C_s5_431));
logic S_s5_432, C_s5_432;
FA FA_s5_432(.A(C_s6_425), .B(C_s6_424), .c_in(C_s6_423), .S(S_s5_432), .c_out(C_s5_432));
logic S_s5_433, C_s5_433;
FA FA_s5_433(.A(C_s6_422), .B(C_s6_421), .c_in(C_s6_420), .S(S_s5_433), .c_out(C_s5_433));
logic S_s5_440, C_s5_440;
FA FA_s5_440(.A(S_s6_445), .B(S_s6_444), .c_in(S_s6_443), .S(S_s5_440), .c_out(C_s5_440));
logic S_s5_441, C_s5_441;
FA FA_s5_441(.A(S_s6_442), .B(S_s6_441), .c_in(S_s6_440), .S(S_s5_441), .c_out(C_s5_441));
logic S_s5_442, C_s5_442;
FA FA_s5_442(.A(C_s6_435), .B(C_s6_434), .c_in(C_s6_433), .S(S_s5_442), .c_out(C_s5_442));
logic S_s5_443, C_s5_443;
FA FA_s5_443(.A(C_s6_432), .B(C_s6_431), .c_in(C_s6_430), .S(S_s5_443), .c_out(C_s5_443));
logic S_s5_450, C_s5_450;
FA FA_s5_450(.A(S_s6_455), .B(S_s6_454), .c_in(S_s6_453), .S(S_s5_450), .c_out(C_s5_450));
logic S_s5_451, C_s5_451;
FA FA_s5_451(.A(S_s6_452), .B(S_s6_451), .c_in(S_s6_450), .S(S_s5_451), .c_out(C_s5_451));
logic S_s5_452, C_s5_452;
FA FA_s5_452(.A(C_s6_445), .B(C_s6_444), .c_in(C_s6_443), .S(S_s5_452), .c_out(C_s5_452));
logic S_s5_453, C_s5_453;
FA FA_s5_453(.A(C_s6_442), .B(C_s6_441), .c_in(C_s6_440), .S(S_s5_453), .c_out(C_s5_453));
logic S_s5_460, C_s5_460;
FA FA_s5_460(.A(S_s6_464), .B(S_s6_463), .c_in(S_s6_462), .S(S_s5_460), .c_out(C_s5_460));
logic S_s5_461, C_s5_461;
FA FA_s5_461(.A(S_s6_461), .B(S_s6_460), .c_in(C_s6_455), .S(S_s5_461), .c_out(C_s5_461));
logic S_s5_462, C_s5_462;
FA FA_s5_462(.A(C_s6_454), .B(C_s6_453), .c_in(C_s6_452), .S(S_s5_462), .c_out(C_s5_462));
logic S_s5_463, C_s5_463;
FA FA_s5_463(.A(C_s6_451), .B(C_s6_450), .c_in(comb[30][16]), .S(S_s5_463), .c_out(C_s5_463));
logic S_s5_470, C_s5_470;
FA FA_s5_470(.A(S_s6_473), .B(S_s6_472), .c_in(S_s6_471), .S(S_s5_470), .c_out(C_s5_470));
logic S_s5_471, C_s5_471;
FA FA_s5_471(.A(S_s6_470), .B(C_s6_464), .c_in(C_s6_463), .S(S_s5_471), .c_out(C_s5_471));
logic S_s5_472, C_s5_472;
FA FA_s5_472(.A(C_s6_462), .B(C_s6_461), .c_in(C_s6_460), .S(S_s5_472), .c_out(C_s5_472));
logic S_s5_473, C_s5_473;
FA FA_s5_473(.A(comb[28][19]), .B(comb[29][18]), .c_in(comb[30][17]), .S(S_s5_473), .c_out(C_s5_473));
logic S_s5_480, C_s5_480;
FA FA_s5_480(.A(S_s6_482), .B(S_s6_481), .c_in(S_s6_480), .S(S_s5_480), .c_out(C_s5_480));
logic S_s5_481, C_s5_481;
FA FA_s5_481(.A(C_s6_473), .B(C_s6_472), .c_in(C_s6_471), .S(S_s5_481), .c_out(C_s5_481));
logic S_s5_482, C_s5_482;
FA FA_s5_482(.A(C_s6_470), .B(comb[26][22]), .c_in(comb[27][21]), .S(S_s5_482), .c_out(C_s5_482));
logic S_s5_483, C_s5_483;
FA FA_s5_483(.A(comb[28][20]), .B(comb[29][19]), .c_in(comb[30][18]), .S(S_s5_483), .c_out(C_s5_483));
logic S_s5_490, C_s5_490;
FA FA_s5_490(.A(S_s6_491), .B(S_s6_490), .c_in(C_s6_482), .S(S_s5_490), .c_out(C_s5_490));
logic S_s5_491, C_s5_491;
FA FA_s5_491(.A(C_s6_481), .B(C_s6_480), .c_in(comb[24][25]), .S(S_s5_491), .c_out(C_s5_491));
logic S_s5_492, C_s5_492;
FA FA_s5_492(.A(comb[25][24]), .B(comb[26][23]), .c_in(comb[27][22]), .S(S_s5_492), .c_out(C_s5_492));
logic S_s5_493, C_s5_493;
FA FA_s5_493(.A(comb[28][21]), .B(comb[29][20]), .c_in(comb[30][19]), .S(S_s5_493), .c_out(C_s5_493));
logic S_s5_500, C_s5_500;
FA FA_s5_500(.A(S_s6_500), .B(C_s6_491), .c_in(C_s6_490), .S(S_s5_500), .c_out(C_s5_500));
logic S_s5_501, C_s5_501;
FA FA_s5_501(.A(comb[22][28]), .B(comb[23][27]), .c_in(comb[24][26]), .S(S_s5_501), .c_out(C_s5_501));
logic S_s5_502, C_s5_502;
FA FA_s5_502(.A(comb[25][25]), .B(comb[26][24]), .c_in(comb[27][23]), .S(S_s5_502), .c_out(C_s5_502));
logic S_s5_503, C_s5_503;
FA FA_s5_503(.A(comb[28][22]), .B(comb[29][21]), .c_in(comb[30][20]), .S(S_s5_503), .c_out(C_s5_503));
logic S_s5_510, C_s5_510;
FA FA_s5_510(.A(C_s6_500), .B(comb[20][31]), .c_in(comb[21][30]), .S(S_s5_510), .c_out(C_s5_510));
logic S_s5_511, C_s5_511;
FA FA_s5_511(.A(comb[22][29]), .B(comb[23][28]), .c_in(comb[24][27]), .S(S_s5_511), .c_out(C_s5_511));
logic S_s5_512, C_s5_512;
FA FA_s5_512(.A(comb[25][26]), .B(comb[26][25]), .c_in(comb[27][24]), .S(S_s5_512), .c_out(C_s5_512));
logic S_s5_513, C_s5_513;
FA FA_s5_513(.A(comb[28][23]), .B(comb[29][22]), .c_in(comb[30][21]), .S(S_s5_513), .c_out(C_s5_513));
logic S_s5_520, C_s5_520;
FA FA_s5_520(.A(comb[21][31]), .B(comb[22][30]), .c_in(comb[23][29]), .S(S_s5_520), .c_out(C_s5_520));
logic S_s5_521, C_s5_521;
FA FA_s5_521(.A(comb[24][28]), .B(comb[25][27]), .c_in(comb[26][26]), .S(S_s5_521), .c_out(C_s5_521));
logic S_s5_522, C_s5_522;
FA FA_s5_522(.A(comb[27][25]), .B(comb[28][24]), .c_in(comb[29][23]), .S(S_s5_522), .c_out(C_s5_522));
logic S_s5_530, C_s5_530;
FA FA_s5_530(.A(comb[22][31]), .B(comb[23][30]), .c_in(comb[24][29]), .S(S_s5_530), .c_out(C_s5_530));
logic S_s5_531, C_s5_531;
FA FA_s5_531(.A(comb[25][28]), .B(comb[26][27]), .c_in(comb[27][26]), .S(S_s5_531), .c_out(C_s5_531));
logic S_s5_540, C_s5_540;
FA FA_s5_540(.A(comb[23][31]), .B(comb[24][30]), .c_in(comb[25][29]), .S(S_s5_540), .c_out(C_s5_540));
// stage 5 end ======================================================================================================= 

// stage 4 begin ======================================================================================================= 
logic S_s4_60, C_s4_60;
HA HA_s4_60(.A(comb[0][6]), .B(comb[1][5]), .S(S_s4_60), .c_out(C_s4_60));
logic S_s4_70, C_s4_70;
FA FA_s4_70(.A(comb[0][7]), .B(comb[1][6]), .c_in(comb[2][5]), .S(S_s4_70), .c_out(C_s4_70));
logic S_s4_71, C_s4_71;
HA HA_s4_71(.A(comb[3][4]), .B(comb[4][3]), .S(S_s4_71), .c_out(C_s4_71));
logic S_s4_80, C_s4_80;
FA FA_s4_80(.A(comb[0][8]), .B(comb[1][7]), .c_in(comb[2][6]), .S(S_s4_80), .c_out(C_s4_80));
logic S_s4_81, C_s4_81;
FA FA_s4_81(.A(comb[3][5]), .B(comb[4][4]), .c_in(comb[5][3]), .S(S_s4_81), .c_out(C_s4_81));
logic S_s4_82, C_s4_82;
HA HA_s4_82(.A(comb[6][2]), .B(comb[7][1]), .S(S_s4_82), .c_out(C_s4_82));
logic S_s4_90, C_s4_90;
FA FA_s4_90(.A(S_s5_90), .B(comb[2][7]), .c_in(comb[3][6]), .S(S_s4_90), .c_out(C_s4_90));
logic S_s4_91, C_s4_91;
FA FA_s4_91(.A(comb[4][5]), .B(comb[5][4]), .c_in(comb[6][3]), .S(S_s4_91), .c_out(C_s4_91));
logic S_s4_92, C_s4_92;
FA FA_s4_92(.A(comb[7][2]), .B(comb[8][1]), .c_in(comb[9][0]), .S(S_s4_92), .c_out(C_s4_92));
logic S_s4_100, C_s4_100;
FA FA_s4_100(.A(S_s5_101), .B(S_s5_100), .c_in(C_s5_90), .S(S_s4_100), .c_out(C_s4_100));
logic S_s4_101, C_s4_101;
FA FA_s4_101(.A(comb[5][5]), .B(comb[6][4]), .c_in(comb[7][3]), .S(S_s4_101), .c_out(C_s4_101));
logic S_s4_102, C_s4_102;
FA FA_s4_102(.A(comb[8][2]), .B(comb[9][1]), .c_in(comb[10][0]), .S(S_s4_102), .c_out(C_s4_102));
logic S_s4_110, C_s4_110;
FA FA_s4_110(.A(S_s5_112), .B(S_s5_111), .c_in(S_s5_110), .S(S_s4_110), .c_out(C_s4_110));
logic S_s4_111, C_s4_111;
FA FA_s4_111(.A(C_s5_101), .B(C_s5_100), .c_in(comb[8][3]), .S(S_s4_111), .c_out(C_s4_111));
logic S_s4_112, C_s4_112;
FA FA_s4_112(.A(comb[9][2]), .B(comb[10][1]), .c_in(comb[11][0]), .S(S_s4_112), .c_out(C_s4_112));
logic S_s4_120, C_s4_120;
FA FA_s4_120(.A(S_s5_123), .B(S_s5_122), .c_in(S_s5_121), .S(S_s4_120), .c_out(C_s4_120));
logic S_s4_121, C_s4_121;
FA FA_s4_121(.A(S_s5_120), .B(C_s5_112), .c_in(C_s5_111), .S(S_s4_121), .c_out(C_s4_121));
logic S_s4_122, C_s4_122;
FA FA_s4_122(.A(C_s5_110), .B(comb[11][1]), .c_in(comb[12][0]), .S(S_s4_122), .c_out(C_s4_122));
logic S_s4_130, C_s4_130;
FA FA_s4_130(.A(S_s5_133), .B(S_s5_132), .c_in(S_s5_131), .S(S_s4_130), .c_out(C_s4_130));
logic S_s4_131, C_s4_131;
FA FA_s4_131(.A(S_s5_130), .B(C_s5_123), .c_in(C_s5_122), .S(S_s4_131), .c_out(C_s4_131));
logic S_s4_132, C_s4_132;
FA FA_s4_132(.A(C_s5_121), .B(C_s5_120), .c_in(comb[13][0]), .S(S_s4_132), .c_out(C_s4_132));
logic S_s4_140, C_s4_140;
FA FA_s4_140(.A(S_s5_143), .B(S_s5_142), .c_in(S_s5_141), .S(S_s4_140), .c_out(C_s4_140));
logic S_s4_141, C_s4_141;
FA FA_s4_141(.A(S_s5_140), .B(C_s5_133), .c_in(C_s5_132), .S(S_s4_141), .c_out(C_s4_141));
logic S_s4_142, C_s4_142;
FA FA_s4_142(.A(C_s5_131), .B(C_s5_130), .c_in(comb[14][0]), .S(S_s4_142), .c_out(C_s4_142));
logic S_s4_150, C_s4_150;
FA FA_s4_150(.A(S_s5_153), .B(S_s5_152), .c_in(S_s5_151), .S(S_s4_150), .c_out(C_s4_150));
logic S_s4_151, C_s4_151;
FA FA_s4_151(.A(S_s5_150), .B(C_s5_143), .c_in(C_s5_142), .S(S_s4_151), .c_out(C_s4_151));
logic S_s4_152, C_s4_152;
FA FA_s4_152(.A(C_s5_141), .B(C_s5_140), .c_in(comb[15][0]), .S(S_s4_152), .c_out(C_s4_152));
logic S_s4_160, C_s4_160;
FA FA_s4_160(.A(S_s5_163), .B(S_s5_162), .c_in(S_s5_161), .S(S_s4_160), .c_out(C_s4_160));
logic S_s4_161, C_s4_161;
FA FA_s4_161(.A(S_s5_160), .B(C_s5_153), .c_in(C_s5_152), .S(S_s4_161), .c_out(C_s4_161));
logic S_s4_162, C_s4_162;
FA FA_s4_162(.A(C_s5_151), .B(C_s5_150), .c_in(comb[16][0]), .S(S_s4_162), .c_out(C_s4_162));
logic S_s4_170, C_s4_170;
FA FA_s4_170(.A(S_s5_173), .B(S_s5_172), .c_in(S_s5_171), .S(S_s4_170), .c_out(C_s4_170));
logic S_s4_171, C_s4_171;
FA FA_s4_171(.A(S_s5_170), .B(C_s5_163), .c_in(C_s5_162), .S(S_s4_171), .c_out(C_s4_171));
logic S_s4_172, C_s4_172;
FA FA_s4_172(.A(C_s5_161), .B(C_s5_160), .c_in(comb[17][0]), .S(S_s4_172), .c_out(C_s4_172));
logic S_s4_180, C_s4_180;
FA FA_s4_180(.A(S_s5_183), .B(S_s5_182), .c_in(S_s5_181), .S(S_s4_180), .c_out(C_s4_180));
logic S_s4_181, C_s4_181;
FA FA_s4_181(.A(S_s5_180), .B(C_s5_173), .c_in(C_s5_172), .S(S_s4_181), .c_out(C_s4_181));
logic S_s4_182, C_s4_182;
FA FA_s4_182(.A(C_s5_171), .B(C_s5_170), .c_in(comb[18][0]), .S(S_s4_182), .c_out(C_s4_182));
logic S_s4_190, C_s4_190;
FA FA_s4_190(.A(S_s5_193), .B(S_s5_192), .c_in(S_s5_191), .S(S_s4_190), .c_out(C_s4_190));
logic S_s4_191, C_s4_191;
FA FA_s4_191(.A(S_s5_190), .B(C_s5_183), .c_in(C_s5_182), .S(S_s4_191), .c_out(C_s4_191));
logic S_s4_192, C_s4_192;
FA FA_s4_192(.A(C_s5_181), .B(C_s5_180), .c_in(comb[19][0]), .S(S_s4_192), .c_out(C_s4_192));
logic S_s4_200, C_s4_200;
FA FA_s4_200(.A(S_s5_203), .B(S_s5_202), .c_in(S_s5_201), .S(S_s4_200), .c_out(C_s4_200));
logic S_s4_201, C_s4_201;
FA FA_s4_201(.A(S_s5_200), .B(C_s5_193), .c_in(C_s5_192), .S(S_s4_201), .c_out(C_s4_201));
logic S_s4_202, C_s4_202;
FA FA_s4_202(.A(C_s5_191), .B(C_s5_190), .c_in(comb[20][0]), .S(S_s4_202), .c_out(C_s4_202));
logic S_s4_210, C_s4_210;
FA FA_s4_210(.A(S_s5_213), .B(S_s5_212), .c_in(S_s5_211), .S(S_s4_210), .c_out(C_s4_210));
logic S_s4_211, C_s4_211;
FA FA_s4_211(.A(S_s5_210), .B(C_s5_203), .c_in(C_s5_202), .S(S_s4_211), .c_out(C_s4_211));
logic S_s4_212, C_s4_212;
FA FA_s4_212(.A(C_s5_201), .B(C_s5_200), .c_in(comb[21][0]), .S(S_s4_212), .c_out(C_s4_212));
logic S_s4_220, C_s4_220;
FA FA_s4_220(.A(S_s5_223), .B(S_s5_222), .c_in(S_s5_221), .S(S_s4_220), .c_out(C_s4_220));
logic S_s4_221, C_s4_221;
FA FA_s4_221(.A(S_s5_220), .B(C_s5_213), .c_in(C_s5_212), .S(S_s4_221), .c_out(C_s4_221));
logic S_s4_222, C_s4_222;
FA FA_s4_222(.A(C_s5_211), .B(C_s5_210), .c_in(comb[22][0]), .S(S_s4_222), .c_out(C_s4_222));
logic S_s4_230, C_s4_230;
FA FA_s4_230(.A(S_s5_233), .B(S_s5_232), .c_in(S_s5_231), .S(S_s4_230), .c_out(C_s4_230));
logic S_s4_231, C_s4_231;
FA FA_s4_231(.A(S_s5_230), .B(C_s5_223), .c_in(C_s5_222), .S(S_s4_231), .c_out(C_s4_231));
logic S_s4_232, C_s4_232;
FA FA_s4_232(.A(C_s5_221), .B(C_s5_220), .c_in(comb[23][0]), .S(S_s4_232), .c_out(C_s4_232));
logic S_s4_240, C_s4_240;
FA FA_s4_240(.A(S_s5_243), .B(S_s5_242), .c_in(S_s5_241), .S(S_s4_240), .c_out(C_s4_240));
logic S_s4_241, C_s4_241;
FA FA_s4_241(.A(S_s5_240), .B(C_s5_233), .c_in(C_s5_232), .S(S_s4_241), .c_out(C_s4_241));
logic S_s4_242, C_s4_242;
FA FA_s4_242(.A(C_s5_231), .B(C_s5_230), .c_in(comb[24][0]), .S(S_s4_242), .c_out(C_s4_242));
logic S_s4_250, C_s4_250;
FA FA_s4_250(.A(S_s5_253), .B(S_s5_252), .c_in(S_s5_251), .S(S_s4_250), .c_out(C_s4_250));
logic S_s4_251, C_s4_251;
FA FA_s4_251(.A(S_s5_250), .B(C_s5_243), .c_in(C_s5_242), .S(S_s4_251), .c_out(C_s4_251));
logic S_s4_252, C_s4_252;
FA FA_s4_252(.A(C_s5_241), .B(C_s5_240), .c_in(comb[25][0]), .S(S_s4_252), .c_out(C_s4_252));
logic S_s4_260, C_s4_260;
FA FA_s4_260(.A(S_s5_263), .B(S_s5_262), .c_in(S_s5_261), .S(S_s4_260), .c_out(C_s4_260));
logic S_s4_261, C_s4_261;
FA FA_s4_261(.A(S_s5_260), .B(C_s5_253), .c_in(C_s5_252), .S(S_s4_261), .c_out(C_s4_261));
logic S_s4_262, C_s4_262;
FA FA_s4_262(.A(C_s5_251), .B(C_s5_250), .c_in(comb[26][0]), .S(S_s4_262), .c_out(C_s4_262));
logic S_s4_270, C_s4_270;
FA FA_s4_270(.A(S_s5_273), .B(S_s5_272), .c_in(S_s5_271), .S(S_s4_270), .c_out(C_s4_270));
logic S_s4_271, C_s4_271;
FA FA_s4_271(.A(S_s5_270), .B(C_s5_263), .c_in(C_s5_262), .S(S_s4_271), .c_out(C_s4_271));
logic S_s4_272, C_s4_272;
FA FA_s4_272(.A(C_s5_261), .B(C_s5_260), .c_in(comb[27][0]), .S(S_s4_272), .c_out(C_s4_272));
logic S_s4_280, C_s4_280;
FA FA_s4_280(.A(S_s5_283), .B(S_s5_282), .c_in(S_s5_281), .S(S_s4_280), .c_out(C_s4_280));
logic S_s4_281, C_s4_281;
FA FA_s4_281(.A(S_s5_280), .B(C_s5_273), .c_in(C_s5_272), .S(S_s4_281), .c_out(C_s4_281));
logic S_s4_282, C_s4_282;
FA FA_s4_282(.A(C_s5_271), .B(C_s5_270), .c_in(comb[28][0]), .S(S_s4_282), .c_out(C_s4_282));
logic S_s4_290, C_s4_290;
FA FA_s4_290(.A(S_s5_293), .B(S_s5_292), .c_in(S_s5_291), .S(S_s4_290), .c_out(C_s4_290));
logic S_s4_291, C_s4_291;
FA FA_s4_291(.A(S_s5_290), .B(C_s5_283), .c_in(C_s5_282), .S(S_s4_291), .c_out(C_s4_291));
logic S_s4_292, C_s4_292;
FA FA_s4_292(.A(C_s5_281), .B(C_s5_280), .c_in(comb[29][0]), .S(S_s4_292), .c_out(C_s4_292));
logic S_s4_300, C_s4_300;
FA FA_s4_300(.A(S_s5_303), .B(S_s5_302), .c_in(S_s5_301), .S(S_s4_300), .c_out(C_s4_300));
logic S_s4_301, C_s4_301;
FA FA_s4_301(.A(S_s5_300), .B(C_s5_293), .c_in(C_s5_292), .S(S_s4_301), .c_out(C_s4_301));
logic S_s4_302, C_s4_302;
FA FA_s4_302(.A(C_s5_291), .B(C_s5_290), .c_in(comb[30][0]), .S(S_s4_302), .c_out(C_s4_302));
logic S_s4_310, C_s4_310;
FA FA_s4_310(.A(S_s5_313), .B(S_s5_312), .c_in(S_s5_311), .S(S_s4_310), .c_out(C_s4_310));
logic S_s4_311, C_s4_311;
FA FA_s4_311(.A(S_s5_310), .B(C_s5_303), .c_in(C_s5_302), .S(S_s4_311), .c_out(C_s4_311));
logic S_s4_312, C_s4_312;
FA FA_s4_312(.A(C_s5_301), .B(C_s5_300), .c_in(comb[31][0]), .S(S_s4_312), .c_out(C_s4_312));
logic S_s4_320, C_s4_320;
FA FA_s4_320(.A(S_s5_323), .B(S_s5_322), .c_in(S_s5_321), .S(S_s4_320), .c_out(C_s4_320));
logic S_s4_321, C_s4_321;
FA FA_s4_321(.A(S_s5_320), .B(C_s5_313), .c_in(C_s5_312), .S(S_s4_321), .c_out(C_s4_321));
logic S_s4_322, C_s4_322;
FA FA_s4_322(.A(C_s5_311), .B(C_s5_310), .c_in(comb[31][1]), .S(S_s4_322), .c_out(C_s4_322));
logic S_s4_330, C_s4_330;
FA FA_s4_330(.A(S_s5_333), .B(S_s5_332), .c_in(S_s5_331), .S(S_s4_330), .c_out(C_s4_330));
logic S_s4_331, C_s4_331;
FA FA_s4_331(.A(S_s5_330), .B(C_s5_323), .c_in(C_s5_322), .S(S_s4_331), .c_out(C_s4_331));
logic S_s4_332, C_s4_332;
FA FA_s4_332(.A(C_s5_321), .B(C_s5_320), .c_in(comb[31][2]), .S(S_s4_332), .c_out(C_s4_332));
logic S_s4_340, C_s4_340;
FA FA_s4_340(.A(S_s5_343), .B(S_s5_342), .c_in(S_s5_341), .S(S_s4_340), .c_out(C_s4_340));
logic S_s4_341, C_s4_341;
FA FA_s4_341(.A(S_s5_340), .B(C_s5_333), .c_in(C_s5_332), .S(S_s4_341), .c_out(C_s4_341));
logic S_s4_342, C_s4_342;
FA FA_s4_342(.A(C_s5_331), .B(C_s5_330), .c_in(comb[31][3]), .S(S_s4_342), .c_out(C_s4_342));
logic S_s4_350, C_s4_350;
FA FA_s4_350(.A(S_s5_353), .B(S_s5_352), .c_in(S_s5_351), .S(S_s4_350), .c_out(C_s4_350));
logic S_s4_351, C_s4_351;
FA FA_s4_351(.A(S_s5_350), .B(C_s5_343), .c_in(C_s5_342), .S(S_s4_351), .c_out(C_s4_351));
logic S_s4_352, C_s4_352;
FA FA_s4_352(.A(C_s5_341), .B(C_s5_340), .c_in(comb[31][4]), .S(S_s4_352), .c_out(C_s4_352));
logic S_s4_360, C_s4_360;
FA FA_s4_360(.A(S_s5_363), .B(S_s5_362), .c_in(S_s5_361), .S(S_s4_360), .c_out(C_s4_360));
logic S_s4_361, C_s4_361;
FA FA_s4_361(.A(S_s5_360), .B(C_s5_353), .c_in(C_s5_352), .S(S_s4_361), .c_out(C_s4_361));
logic S_s4_362, C_s4_362;
FA FA_s4_362(.A(C_s5_351), .B(C_s5_350), .c_in(comb[31][5]), .S(S_s4_362), .c_out(C_s4_362));
logic S_s4_370, C_s4_370;
FA FA_s4_370(.A(S_s5_373), .B(S_s5_372), .c_in(S_s5_371), .S(S_s4_370), .c_out(C_s4_370));
logic S_s4_371, C_s4_371;
FA FA_s4_371(.A(S_s5_370), .B(C_s5_363), .c_in(C_s5_362), .S(S_s4_371), .c_out(C_s4_371));
logic S_s4_372, C_s4_372;
FA FA_s4_372(.A(C_s5_361), .B(C_s5_360), .c_in(comb[31][6]), .S(S_s4_372), .c_out(C_s4_372));
logic S_s4_380, C_s4_380;
FA FA_s4_380(.A(S_s5_383), .B(S_s5_382), .c_in(S_s5_381), .S(S_s4_380), .c_out(C_s4_380));
logic S_s4_381, C_s4_381;
FA FA_s4_381(.A(S_s5_380), .B(C_s5_373), .c_in(C_s5_372), .S(S_s4_381), .c_out(C_s4_381));
logic S_s4_382, C_s4_382;
FA FA_s4_382(.A(C_s5_371), .B(C_s5_370), .c_in(comb[31][7]), .S(S_s4_382), .c_out(C_s4_382));
logic S_s4_390, C_s4_390;
FA FA_s4_390(.A(S_s5_393), .B(S_s5_392), .c_in(S_s5_391), .S(S_s4_390), .c_out(C_s4_390));
logic S_s4_391, C_s4_391;
FA FA_s4_391(.A(S_s5_390), .B(C_s5_383), .c_in(C_s5_382), .S(S_s4_391), .c_out(C_s4_391));
logic S_s4_392, C_s4_392;
FA FA_s4_392(.A(C_s5_381), .B(C_s5_380), .c_in(comb[31][8]), .S(S_s4_392), .c_out(C_s4_392));
logic S_s4_400, C_s4_400;
FA FA_s4_400(.A(S_s5_403), .B(S_s5_402), .c_in(S_s5_401), .S(S_s4_400), .c_out(C_s4_400));
logic S_s4_401, C_s4_401;
FA FA_s4_401(.A(S_s5_400), .B(C_s5_393), .c_in(C_s5_392), .S(S_s4_401), .c_out(C_s4_401));
logic S_s4_402, C_s4_402;
FA FA_s4_402(.A(C_s5_391), .B(C_s5_390), .c_in(comb[31][9]), .S(S_s4_402), .c_out(C_s4_402));
logic S_s4_410, C_s4_410;
FA FA_s4_410(.A(S_s5_413), .B(S_s5_412), .c_in(S_s5_411), .S(S_s4_410), .c_out(C_s4_410));
logic S_s4_411, C_s4_411;
FA FA_s4_411(.A(S_s5_410), .B(C_s5_403), .c_in(C_s5_402), .S(S_s4_411), .c_out(C_s4_411));
logic S_s4_412, C_s4_412;
FA FA_s4_412(.A(C_s5_401), .B(C_s5_400), .c_in(comb[31][10]), .S(S_s4_412), .c_out(C_s4_412));
logic S_s4_420, C_s4_420;
FA FA_s4_420(.A(S_s5_423), .B(S_s5_422), .c_in(S_s5_421), .S(S_s4_420), .c_out(C_s4_420));
logic S_s4_421, C_s4_421;
FA FA_s4_421(.A(S_s5_420), .B(C_s5_413), .c_in(C_s5_412), .S(S_s4_421), .c_out(C_s4_421));
logic S_s4_422, C_s4_422;
FA FA_s4_422(.A(C_s5_411), .B(C_s5_410), .c_in(comb[31][11]), .S(S_s4_422), .c_out(C_s4_422));
logic S_s4_430, C_s4_430;
FA FA_s4_430(.A(S_s5_433), .B(S_s5_432), .c_in(S_s5_431), .S(S_s4_430), .c_out(C_s4_430));
logic S_s4_431, C_s4_431;
FA FA_s4_431(.A(S_s5_430), .B(C_s5_423), .c_in(C_s5_422), .S(S_s4_431), .c_out(C_s4_431));
logic S_s4_432, C_s4_432;
FA FA_s4_432(.A(C_s5_421), .B(C_s5_420), .c_in(comb[31][12]), .S(S_s4_432), .c_out(C_s4_432));
logic S_s4_440, C_s4_440;
FA FA_s4_440(.A(S_s5_443), .B(S_s5_442), .c_in(S_s5_441), .S(S_s4_440), .c_out(C_s4_440));
logic S_s4_441, C_s4_441;
FA FA_s4_441(.A(S_s5_440), .B(C_s5_433), .c_in(C_s5_432), .S(S_s4_441), .c_out(C_s4_441));
logic S_s4_442, C_s4_442;
FA FA_s4_442(.A(C_s5_431), .B(C_s5_430), .c_in(comb[31][13]), .S(S_s4_442), .c_out(C_s4_442));
logic S_s4_450, C_s4_450;
FA FA_s4_450(.A(S_s5_453), .B(S_s5_452), .c_in(S_s5_451), .S(S_s4_450), .c_out(C_s4_450));
logic S_s4_451, C_s4_451;
FA FA_s4_451(.A(S_s5_450), .B(C_s5_443), .c_in(C_s5_442), .S(S_s4_451), .c_out(C_s4_451));
logic S_s4_452, C_s4_452;
FA FA_s4_452(.A(C_s5_441), .B(C_s5_440), .c_in(comb[31][14]), .S(S_s4_452), .c_out(C_s4_452));
logic S_s4_460, C_s4_460;
FA FA_s4_460(.A(S_s5_463), .B(S_s5_462), .c_in(S_s5_461), .S(S_s4_460), .c_out(C_s4_460));
logic S_s4_461, C_s4_461;
FA FA_s4_461(.A(S_s5_460), .B(C_s5_453), .c_in(C_s5_452), .S(S_s4_461), .c_out(C_s4_461));
logic S_s4_462, C_s4_462;
FA FA_s4_462(.A(C_s5_451), .B(C_s5_450), .c_in(comb[31][15]), .S(S_s4_462), .c_out(C_s4_462));
logic S_s4_470, C_s4_470;
FA FA_s4_470(.A(S_s5_473), .B(S_s5_472), .c_in(S_s5_471), .S(S_s4_470), .c_out(C_s4_470));
logic S_s4_471, C_s4_471;
FA FA_s4_471(.A(S_s5_470), .B(C_s5_463), .c_in(C_s5_462), .S(S_s4_471), .c_out(C_s4_471));
logic S_s4_472, C_s4_472;
FA FA_s4_472(.A(C_s5_461), .B(C_s5_460), .c_in(comb[31][16]), .S(S_s4_472), .c_out(C_s4_472));
logic S_s4_480, C_s4_480;
FA FA_s4_480(.A(S_s5_483), .B(S_s5_482), .c_in(S_s5_481), .S(S_s4_480), .c_out(C_s4_480));
logic S_s4_481, C_s4_481;
FA FA_s4_481(.A(S_s5_480), .B(C_s5_473), .c_in(C_s5_472), .S(S_s4_481), .c_out(C_s4_481));
logic S_s4_482, C_s4_482;
FA FA_s4_482(.A(C_s5_471), .B(C_s5_470), .c_in(comb[31][17]), .S(S_s4_482), .c_out(C_s4_482));
logic S_s4_490, C_s4_490;
FA FA_s4_490(.A(S_s5_493), .B(S_s5_492), .c_in(S_s5_491), .S(S_s4_490), .c_out(C_s4_490));
logic S_s4_491, C_s4_491;
FA FA_s4_491(.A(S_s5_490), .B(C_s5_483), .c_in(C_s5_482), .S(S_s4_491), .c_out(C_s4_491));
logic S_s4_492, C_s4_492;
FA FA_s4_492(.A(C_s5_481), .B(C_s5_480), .c_in(comb[31][18]), .S(S_s4_492), .c_out(C_s4_492));
logic S_s4_500, C_s4_500;
FA FA_s4_500(.A(S_s5_503), .B(S_s5_502), .c_in(S_s5_501), .S(S_s4_500), .c_out(C_s4_500));
logic S_s4_501, C_s4_501;
FA FA_s4_501(.A(S_s5_500), .B(C_s5_493), .c_in(C_s5_492), .S(S_s4_501), .c_out(C_s4_501));
logic S_s4_502, C_s4_502;
FA FA_s4_502(.A(C_s5_491), .B(C_s5_490), .c_in(comb[31][19]), .S(S_s4_502), .c_out(C_s4_502));
logic S_s4_510, C_s4_510;
FA FA_s4_510(.A(S_s5_513), .B(S_s5_512), .c_in(S_s5_511), .S(S_s4_510), .c_out(C_s4_510));
logic S_s4_511, C_s4_511;
FA FA_s4_511(.A(S_s5_510), .B(C_s5_503), .c_in(C_s5_502), .S(S_s4_511), .c_out(C_s4_511));
logic S_s4_512, C_s4_512;
FA FA_s4_512(.A(C_s5_501), .B(C_s5_500), .c_in(comb[31][20]), .S(S_s4_512), .c_out(C_s4_512));
logic S_s4_520, C_s4_520;
FA FA_s4_520(.A(S_s5_522), .B(S_s5_521), .c_in(S_s5_520), .S(S_s4_520), .c_out(C_s4_520));
logic S_s4_521, C_s4_521;
FA FA_s4_521(.A(C_s5_513), .B(C_s5_512), .c_in(C_s5_511), .S(S_s4_521), .c_out(C_s4_521));
logic S_s4_522, C_s4_522;
FA FA_s4_522(.A(C_s5_510), .B(comb[30][22]), .c_in(comb[31][21]), .S(S_s4_522), .c_out(C_s4_522));
logic S_s4_530, C_s4_530;
FA FA_s4_530(.A(S_s5_531), .B(S_s5_530), .c_in(C_s5_522), .S(S_s4_530), .c_out(C_s4_530));
logic S_s4_531, C_s4_531;
FA FA_s4_531(.A(C_s5_521), .B(C_s5_520), .c_in(comb[28][25]), .S(S_s4_531), .c_out(C_s4_531));
logic S_s4_532, C_s4_532;
FA FA_s4_532(.A(comb[29][24]), .B(comb[30][23]), .c_in(comb[31][22]), .S(S_s4_532), .c_out(C_s4_532));
logic S_s4_540, C_s4_540;
FA FA_s4_540(.A(S_s5_540), .B(C_s5_531), .c_in(C_s5_530), .S(S_s4_540), .c_out(C_s4_540));
logic S_s4_541, C_s4_541;
FA FA_s4_541(.A(comb[26][28]), .B(comb[27][27]), .c_in(comb[28][26]), .S(S_s4_541), .c_out(C_s4_541));
logic S_s4_542, C_s4_542;
FA FA_s4_542(.A(comb[29][25]), .B(comb[30][24]), .c_in(comb[31][23]), .S(S_s4_542), .c_out(C_s4_542));
logic S_s4_550, C_s4_550;
FA FA_s4_550(.A(C_s5_540), .B(comb[24][31]), .c_in(comb[25][30]), .S(S_s4_550), .c_out(C_s4_550));
logic S_s4_551, C_s4_551;
FA FA_s4_551(.A(comb[26][29]), .B(comb[27][28]), .c_in(comb[28][27]), .S(S_s4_551), .c_out(C_s4_551));
logic S_s4_552, C_s4_552;
FA FA_s4_552(.A(comb[29][26]), .B(comb[30][25]), .c_in(comb[31][24]), .S(S_s4_552), .c_out(C_s4_552));
logic S_s4_560, C_s4_560;
FA FA_s4_560(.A(comb[25][31]), .B(comb[26][30]), .c_in(comb[27][29]), .S(S_s4_560), .c_out(C_s4_560));
logic S_s4_561, C_s4_561;
FA FA_s4_561(.A(comb[28][28]), .B(comb[29][27]), .c_in(comb[30][26]), .S(S_s4_561), .c_out(C_s4_561));
logic S_s4_570, C_s4_570;
FA FA_s4_570(.A(comb[26][31]), .B(comb[27][30]), .c_in(comb[28][29]), .S(S_s4_570), .c_out(C_s4_570));
// stage 4 end ======================================================================================================= 

// stage 3 begin ======================================================================================================= 
logic S_s3_40, C_s3_40;
HA HA_s3_40(.A(comb[0][4]), .B(comb[1][3]), .S(S_s3_40), .c_out(C_s3_40));
logic S_s3_50, C_s3_50;
FA FA_s3_50(.A(comb[0][5]), .B(comb[1][4]), .c_in(comb[2][3]), .S(S_s3_50), .c_out(C_s3_50));
logic S_s3_51, C_s3_51;
HA HA_s3_51(.A(comb[3][2]), .B(comb[4][1]), .S(S_s3_51), .c_out(C_s3_51));
logic S_s3_60, C_s3_60;
FA FA_s3_60(.A(S_s4_60), .B(comb[2][4]), .c_in(comb[3][3]), .S(S_s3_60), .c_out(C_s3_60));
logic S_s3_61, C_s3_61;
FA FA_s3_61(.A(comb[4][2]), .B(comb[5][1]), .c_in(comb[6][0]), .S(S_s3_61), .c_out(C_s3_61));
logic S_s3_70, C_s3_70;
FA FA_s3_70(.A(S_s4_71), .B(S_s4_70), .c_in(C_s4_60), .S(S_s3_70), .c_out(C_s3_70));
logic S_s3_71, C_s3_71;
FA FA_s3_71(.A(comb[5][2]), .B(comb[6][1]), .c_in(comb[7][0]), .S(S_s3_71), .c_out(C_s3_71));
logic S_s3_80, C_s3_80;
FA FA_s3_80(.A(S_s4_82), .B(S_s4_81), .c_in(S_s4_80), .S(S_s3_80), .c_out(C_s3_80));
logic S_s3_81, C_s3_81;
FA FA_s3_81(.A(C_s4_71), .B(C_s4_70), .c_in(comb[8][0]), .S(S_s3_81), .c_out(C_s3_81));
logic S_s3_90, C_s3_90;
FA FA_s3_90(.A(S_s4_92), .B(S_s4_91), .c_in(S_s4_90), .S(S_s3_90), .c_out(C_s3_90));
logic S_s3_91, C_s3_91;
FA FA_s3_91(.A(C_s4_82), .B(C_s4_81), .c_in(C_s4_80), .S(S_s3_91), .c_out(C_s3_91));
logic S_s3_100, C_s3_100;
FA FA_s3_100(.A(S_s4_102), .B(S_s4_101), .c_in(S_s4_100), .S(S_s3_100), .c_out(C_s3_100));
logic S_s3_101, C_s3_101;
FA FA_s3_101(.A(C_s4_92), .B(C_s4_91), .c_in(C_s4_90), .S(S_s3_101), .c_out(C_s3_101));
logic S_s3_110, C_s3_110;
FA FA_s3_110(.A(S_s4_112), .B(S_s4_111), .c_in(S_s4_110), .S(S_s3_110), .c_out(C_s3_110));
logic S_s3_111, C_s3_111;
FA FA_s3_111(.A(C_s4_102), .B(C_s4_101), .c_in(C_s4_100), .S(S_s3_111), .c_out(C_s3_111));
logic S_s3_120, C_s3_120;
FA FA_s3_120(.A(S_s4_122), .B(S_s4_121), .c_in(S_s4_120), .S(S_s3_120), .c_out(C_s3_120));
logic S_s3_121, C_s3_121;
FA FA_s3_121(.A(C_s4_112), .B(C_s4_111), .c_in(C_s4_110), .S(S_s3_121), .c_out(C_s3_121));
logic S_s3_130, C_s3_130;
FA FA_s3_130(.A(S_s4_132), .B(S_s4_131), .c_in(S_s4_130), .S(S_s3_130), .c_out(C_s3_130));
logic S_s3_131, C_s3_131;
FA FA_s3_131(.A(C_s4_122), .B(C_s4_121), .c_in(C_s4_120), .S(S_s3_131), .c_out(C_s3_131));
logic S_s3_140, C_s3_140;
FA FA_s3_140(.A(S_s4_142), .B(S_s4_141), .c_in(S_s4_140), .S(S_s3_140), .c_out(C_s3_140));
logic S_s3_141, C_s3_141;
FA FA_s3_141(.A(C_s4_132), .B(C_s4_131), .c_in(C_s4_130), .S(S_s3_141), .c_out(C_s3_141));
logic S_s3_150, C_s3_150;
FA FA_s3_150(.A(S_s4_152), .B(S_s4_151), .c_in(S_s4_150), .S(S_s3_150), .c_out(C_s3_150));
logic S_s3_151, C_s3_151;
FA FA_s3_151(.A(C_s4_142), .B(C_s4_141), .c_in(C_s4_140), .S(S_s3_151), .c_out(C_s3_151));
logic S_s3_160, C_s3_160;
FA FA_s3_160(.A(S_s4_162), .B(S_s4_161), .c_in(S_s4_160), .S(S_s3_160), .c_out(C_s3_160));
logic S_s3_161, C_s3_161;
FA FA_s3_161(.A(C_s4_152), .B(C_s4_151), .c_in(C_s4_150), .S(S_s3_161), .c_out(C_s3_161));
logic S_s3_170, C_s3_170;
FA FA_s3_170(.A(S_s4_172), .B(S_s4_171), .c_in(S_s4_170), .S(S_s3_170), .c_out(C_s3_170));
logic S_s3_171, C_s3_171;
FA FA_s3_171(.A(C_s4_162), .B(C_s4_161), .c_in(C_s4_160), .S(S_s3_171), .c_out(C_s3_171));
logic S_s3_180, C_s3_180;
FA FA_s3_180(.A(S_s4_182), .B(S_s4_181), .c_in(S_s4_180), .S(S_s3_180), .c_out(C_s3_180));
logic S_s3_181, C_s3_181;
FA FA_s3_181(.A(C_s4_172), .B(C_s4_171), .c_in(C_s4_170), .S(S_s3_181), .c_out(C_s3_181));
logic S_s3_190, C_s3_190;
FA FA_s3_190(.A(S_s4_192), .B(S_s4_191), .c_in(S_s4_190), .S(S_s3_190), .c_out(C_s3_190));
logic S_s3_191, C_s3_191;
FA FA_s3_191(.A(C_s4_182), .B(C_s4_181), .c_in(C_s4_180), .S(S_s3_191), .c_out(C_s3_191));
logic S_s3_200, C_s3_200;
FA FA_s3_200(.A(S_s4_202), .B(S_s4_201), .c_in(S_s4_200), .S(S_s3_200), .c_out(C_s3_200));
logic S_s3_201, C_s3_201;
FA FA_s3_201(.A(C_s4_192), .B(C_s4_191), .c_in(C_s4_190), .S(S_s3_201), .c_out(C_s3_201));
logic S_s3_210, C_s3_210;
FA FA_s3_210(.A(S_s4_212), .B(S_s4_211), .c_in(S_s4_210), .S(S_s3_210), .c_out(C_s3_210));
logic S_s3_211, C_s3_211;
FA FA_s3_211(.A(C_s4_202), .B(C_s4_201), .c_in(C_s4_200), .S(S_s3_211), .c_out(C_s3_211));
logic S_s3_220, C_s3_220;
FA FA_s3_220(.A(S_s4_222), .B(S_s4_221), .c_in(S_s4_220), .S(S_s3_220), .c_out(C_s3_220));
logic S_s3_221, C_s3_221;
FA FA_s3_221(.A(C_s4_212), .B(C_s4_211), .c_in(C_s4_210), .S(S_s3_221), .c_out(C_s3_221));
logic S_s3_230, C_s3_230;
FA FA_s3_230(.A(S_s4_232), .B(S_s4_231), .c_in(S_s4_230), .S(S_s3_230), .c_out(C_s3_230));
logic S_s3_231, C_s3_231;
FA FA_s3_231(.A(C_s4_222), .B(C_s4_221), .c_in(C_s4_220), .S(S_s3_231), .c_out(C_s3_231));
logic S_s3_240, C_s3_240;
FA FA_s3_240(.A(S_s4_242), .B(S_s4_241), .c_in(S_s4_240), .S(S_s3_240), .c_out(C_s3_240));
logic S_s3_241, C_s3_241;
FA FA_s3_241(.A(C_s4_232), .B(C_s4_231), .c_in(C_s4_230), .S(S_s3_241), .c_out(C_s3_241));
logic S_s3_250, C_s3_250;
FA FA_s3_250(.A(S_s4_252), .B(S_s4_251), .c_in(S_s4_250), .S(S_s3_250), .c_out(C_s3_250));
logic S_s3_251, C_s3_251;
FA FA_s3_251(.A(C_s4_242), .B(C_s4_241), .c_in(C_s4_240), .S(S_s3_251), .c_out(C_s3_251));
logic S_s3_260, C_s3_260;
FA FA_s3_260(.A(S_s4_262), .B(S_s4_261), .c_in(S_s4_260), .S(S_s3_260), .c_out(C_s3_260));
logic S_s3_261, C_s3_261;
FA FA_s3_261(.A(C_s4_252), .B(C_s4_251), .c_in(C_s4_250), .S(S_s3_261), .c_out(C_s3_261));
logic S_s3_270, C_s3_270;
FA FA_s3_270(.A(S_s4_272), .B(S_s4_271), .c_in(S_s4_270), .S(S_s3_270), .c_out(C_s3_270));
logic S_s3_271, C_s3_271;
FA FA_s3_271(.A(C_s4_262), .B(C_s4_261), .c_in(C_s4_260), .S(S_s3_271), .c_out(C_s3_271));
logic S_s3_280, C_s3_280;
FA FA_s3_280(.A(S_s4_282), .B(S_s4_281), .c_in(S_s4_280), .S(S_s3_280), .c_out(C_s3_280));
logic S_s3_281, C_s3_281;
FA FA_s3_281(.A(C_s4_272), .B(C_s4_271), .c_in(C_s4_270), .S(S_s3_281), .c_out(C_s3_281));
logic S_s3_290, C_s3_290;
FA FA_s3_290(.A(S_s4_292), .B(S_s4_291), .c_in(S_s4_290), .S(S_s3_290), .c_out(C_s3_290));
logic S_s3_291, C_s3_291;
FA FA_s3_291(.A(C_s4_282), .B(C_s4_281), .c_in(C_s4_280), .S(S_s3_291), .c_out(C_s3_291));
logic S_s3_300, C_s3_300;
FA FA_s3_300(.A(S_s4_302), .B(S_s4_301), .c_in(S_s4_300), .S(S_s3_300), .c_out(C_s3_300));
logic S_s3_301, C_s3_301;
FA FA_s3_301(.A(C_s4_292), .B(C_s4_291), .c_in(C_s4_290), .S(S_s3_301), .c_out(C_s3_301));
logic S_s3_310, C_s3_310;
FA FA_s3_310(.A(S_s4_312), .B(S_s4_311), .c_in(S_s4_310), .S(S_s3_310), .c_out(C_s3_310));
logic S_s3_311, C_s3_311;
FA FA_s3_311(.A(C_s4_302), .B(C_s4_301), .c_in(C_s4_300), .S(S_s3_311), .c_out(C_s3_311));
logic S_s3_320, C_s3_320;
FA FA_s3_320(.A(S_s4_322), .B(S_s4_321), .c_in(S_s4_320), .S(S_s3_320), .c_out(C_s3_320));
logic S_s3_321, C_s3_321;
FA FA_s3_321(.A(C_s4_312), .B(C_s4_311), .c_in(C_s4_310), .S(S_s3_321), .c_out(C_s3_321));
logic S_s3_330, C_s3_330;
FA FA_s3_330(.A(S_s4_332), .B(S_s4_331), .c_in(S_s4_330), .S(S_s3_330), .c_out(C_s3_330));
logic S_s3_331, C_s3_331;
FA FA_s3_331(.A(C_s4_322), .B(C_s4_321), .c_in(C_s4_320), .S(S_s3_331), .c_out(C_s3_331));
logic S_s3_340, C_s3_340;
FA FA_s3_340(.A(S_s4_342), .B(S_s4_341), .c_in(S_s4_340), .S(S_s3_340), .c_out(C_s3_340));
logic S_s3_341, C_s3_341;
FA FA_s3_341(.A(C_s4_332), .B(C_s4_331), .c_in(C_s4_330), .S(S_s3_341), .c_out(C_s3_341));
logic S_s3_350, C_s3_350;
FA FA_s3_350(.A(S_s4_352), .B(S_s4_351), .c_in(S_s4_350), .S(S_s3_350), .c_out(C_s3_350));
logic S_s3_351, C_s3_351;
FA FA_s3_351(.A(C_s4_342), .B(C_s4_341), .c_in(C_s4_340), .S(S_s3_351), .c_out(C_s3_351));
logic S_s3_360, C_s3_360;
FA FA_s3_360(.A(S_s4_362), .B(S_s4_361), .c_in(S_s4_360), .S(S_s3_360), .c_out(C_s3_360));
logic S_s3_361, C_s3_361;
FA FA_s3_361(.A(C_s4_352), .B(C_s4_351), .c_in(C_s4_350), .S(S_s3_361), .c_out(C_s3_361));
logic S_s3_370, C_s3_370;
FA FA_s3_370(.A(S_s4_372), .B(S_s4_371), .c_in(S_s4_370), .S(S_s3_370), .c_out(C_s3_370));
logic S_s3_371, C_s3_371;
FA FA_s3_371(.A(C_s4_362), .B(C_s4_361), .c_in(C_s4_360), .S(S_s3_371), .c_out(C_s3_371));
logic S_s3_380, C_s3_380;
FA FA_s3_380(.A(S_s4_382), .B(S_s4_381), .c_in(S_s4_380), .S(S_s3_380), .c_out(C_s3_380));
logic S_s3_381, C_s3_381;
FA FA_s3_381(.A(C_s4_372), .B(C_s4_371), .c_in(C_s4_370), .S(S_s3_381), .c_out(C_s3_381));
logic S_s3_390, C_s3_390;
FA FA_s3_390(.A(S_s4_392), .B(S_s4_391), .c_in(S_s4_390), .S(S_s3_390), .c_out(C_s3_390));
logic S_s3_391, C_s3_391;
FA FA_s3_391(.A(C_s4_382), .B(C_s4_381), .c_in(C_s4_380), .S(S_s3_391), .c_out(C_s3_391));
logic S_s3_400, C_s3_400;
FA FA_s3_400(.A(S_s4_402), .B(S_s4_401), .c_in(S_s4_400), .S(S_s3_400), .c_out(C_s3_400));
logic S_s3_401, C_s3_401;
FA FA_s3_401(.A(C_s4_392), .B(C_s4_391), .c_in(C_s4_390), .S(S_s3_401), .c_out(C_s3_401));
logic S_s3_410, C_s3_410;
FA FA_s3_410(.A(S_s4_412), .B(S_s4_411), .c_in(S_s4_410), .S(S_s3_410), .c_out(C_s3_410));
logic S_s3_411, C_s3_411;
FA FA_s3_411(.A(C_s4_402), .B(C_s4_401), .c_in(C_s4_400), .S(S_s3_411), .c_out(C_s3_411));
logic S_s3_420, C_s3_420;
FA FA_s3_420(.A(S_s4_422), .B(S_s4_421), .c_in(S_s4_420), .S(S_s3_420), .c_out(C_s3_420));
logic S_s3_421, C_s3_421;
FA FA_s3_421(.A(C_s4_412), .B(C_s4_411), .c_in(C_s4_410), .S(S_s3_421), .c_out(C_s3_421));
logic S_s3_430, C_s3_430;
FA FA_s3_430(.A(S_s4_432), .B(S_s4_431), .c_in(S_s4_430), .S(S_s3_430), .c_out(C_s3_430));
logic S_s3_431, C_s3_431;
FA FA_s3_431(.A(C_s4_422), .B(C_s4_421), .c_in(C_s4_420), .S(S_s3_431), .c_out(C_s3_431));
logic S_s3_440, C_s3_440;
FA FA_s3_440(.A(S_s4_442), .B(S_s4_441), .c_in(S_s4_440), .S(S_s3_440), .c_out(C_s3_440));
logic S_s3_441, C_s3_441;
FA FA_s3_441(.A(C_s4_432), .B(C_s4_431), .c_in(C_s4_430), .S(S_s3_441), .c_out(C_s3_441));
logic S_s3_450, C_s3_450;
FA FA_s3_450(.A(S_s4_452), .B(S_s4_451), .c_in(S_s4_450), .S(S_s3_450), .c_out(C_s3_450));
logic S_s3_451, C_s3_451;
FA FA_s3_451(.A(C_s4_442), .B(C_s4_441), .c_in(C_s4_440), .S(S_s3_451), .c_out(C_s3_451));
logic S_s3_460, C_s3_460;
FA FA_s3_460(.A(S_s4_462), .B(S_s4_461), .c_in(S_s4_460), .S(S_s3_460), .c_out(C_s3_460));
logic S_s3_461, C_s3_461;
FA FA_s3_461(.A(C_s4_452), .B(C_s4_451), .c_in(C_s4_450), .S(S_s3_461), .c_out(C_s3_461));
logic S_s3_470, C_s3_470;
FA FA_s3_470(.A(S_s4_472), .B(S_s4_471), .c_in(S_s4_470), .S(S_s3_470), .c_out(C_s3_470));
logic S_s3_471, C_s3_471;
FA FA_s3_471(.A(C_s4_462), .B(C_s4_461), .c_in(C_s4_460), .S(S_s3_471), .c_out(C_s3_471));
logic S_s3_480, C_s3_480;
FA FA_s3_480(.A(S_s4_482), .B(S_s4_481), .c_in(S_s4_480), .S(S_s3_480), .c_out(C_s3_480));
logic S_s3_481, C_s3_481;
FA FA_s3_481(.A(C_s4_472), .B(C_s4_471), .c_in(C_s4_470), .S(S_s3_481), .c_out(C_s3_481));
logic S_s3_490, C_s3_490;
FA FA_s3_490(.A(S_s4_492), .B(S_s4_491), .c_in(S_s4_490), .S(S_s3_490), .c_out(C_s3_490));
logic S_s3_491, C_s3_491;
FA FA_s3_491(.A(C_s4_482), .B(C_s4_481), .c_in(C_s4_480), .S(S_s3_491), .c_out(C_s3_491));
logic S_s3_500, C_s3_500;
FA FA_s3_500(.A(S_s4_502), .B(S_s4_501), .c_in(S_s4_500), .S(S_s3_500), .c_out(C_s3_500));
logic S_s3_501, C_s3_501;
FA FA_s3_501(.A(C_s4_492), .B(C_s4_491), .c_in(C_s4_490), .S(S_s3_501), .c_out(C_s3_501));
logic S_s3_510, C_s3_510;
FA FA_s3_510(.A(S_s4_512), .B(S_s4_511), .c_in(S_s4_510), .S(S_s3_510), .c_out(C_s3_510));
logic S_s3_511, C_s3_511;
FA FA_s3_511(.A(C_s4_502), .B(C_s4_501), .c_in(C_s4_500), .S(S_s3_511), .c_out(C_s3_511));
logic S_s3_520, C_s3_520;
FA FA_s3_520(.A(S_s4_522), .B(S_s4_521), .c_in(S_s4_520), .S(S_s3_520), .c_out(C_s3_520));
logic S_s3_521, C_s3_521;
FA FA_s3_521(.A(C_s4_512), .B(C_s4_511), .c_in(C_s4_510), .S(S_s3_521), .c_out(C_s3_521));
logic S_s3_530, C_s3_530;
FA FA_s3_530(.A(S_s4_532), .B(S_s4_531), .c_in(S_s4_530), .S(S_s3_530), .c_out(C_s3_530));
logic S_s3_531, C_s3_531;
FA FA_s3_531(.A(C_s4_522), .B(C_s4_521), .c_in(C_s4_520), .S(S_s3_531), .c_out(C_s3_531));
logic S_s3_540, C_s3_540;
FA FA_s3_540(.A(S_s4_542), .B(S_s4_541), .c_in(S_s4_540), .S(S_s3_540), .c_out(C_s3_540));
logic S_s3_541, C_s3_541;
FA FA_s3_541(.A(C_s4_532), .B(C_s4_531), .c_in(C_s4_530), .S(S_s3_541), .c_out(C_s3_541));
logic S_s3_550, C_s3_550;
FA FA_s3_550(.A(S_s4_552), .B(S_s4_551), .c_in(S_s4_550), .S(S_s3_550), .c_out(C_s3_550));
logic S_s3_551, C_s3_551;
FA FA_s3_551(.A(C_s4_542), .B(C_s4_541), .c_in(C_s4_540), .S(S_s3_551), .c_out(C_s3_551));
logic S_s3_560, C_s3_560;
FA FA_s3_560(.A(S_s4_561), .B(S_s4_560), .c_in(C_s4_552), .S(S_s3_560), .c_out(C_s3_560));
logic S_s3_561, C_s3_561;
FA FA_s3_561(.A(C_s4_551), .B(C_s4_550), .c_in(comb[31][25]), .S(S_s3_561), .c_out(C_s3_561));
logic S_s3_570, C_s3_570;
FA FA_s3_570(.A(S_s4_570), .B(C_s4_561), .c_in(C_s4_560), .S(S_s3_570), .c_out(C_s3_570));
logic S_s3_571, C_s3_571;
FA FA_s3_571(.A(comb[29][28]), .B(comb[30][27]), .c_in(comb[31][26]), .S(S_s3_571), .c_out(C_s3_571));
logic S_s3_580, C_s3_580;
FA FA_s3_580(.A(C_s4_570), .B(comb[27][31]), .c_in(comb[28][30]), .S(S_s3_580), .c_out(C_s3_580));
logic S_s3_581, C_s3_581;
FA FA_s3_581(.A(comb[29][29]), .B(comb[30][28]), .c_in(comb[31][27]), .S(S_s3_581), .c_out(C_s3_581));
logic S_s3_590, C_s3_590;
FA FA_s3_590(.A(comb[28][31]), .B(comb[29][30]), .c_in(comb[30][29]), .S(S_s3_590), .c_out(C_s3_590));
// stage 3 end ======================================================================================================= 

// stage 2 begin ======================================================================================================= 
logic S_s2_30, C_s2_30;
HA HA_s2_30(.A(comb[0][3]), .B(comb[1][2]), .S(S_s2_30), .c_out(C_s2_30));
logic S_s2_40, C_s2_40;
FA FA_s2_40(.A(S_s3_40), .B(comb[2][2]), .c_in(comb[3][1]), .S(S_s2_40), .c_out(C_s2_40));
logic S_s2_50, C_s2_50;
FA FA_s2_50(.A(S_s3_51), .B(S_s3_50), .c_in(C_s3_40), .S(S_s2_50), .c_out(C_s2_50));
logic S_s2_60, C_s2_60;
FA FA_s2_60(.A(S_s3_61), .B(S_s3_60), .c_in(C_s3_51), .S(S_s2_60), .c_out(C_s2_60));
logic S_s2_70, C_s2_70;
FA FA_s2_70(.A(S_s3_71), .B(S_s3_70), .c_in(C_s3_61), .S(S_s2_70), .c_out(C_s2_70));
logic S_s2_80, C_s2_80;
FA FA_s2_80(.A(S_s3_81), .B(S_s3_80), .c_in(C_s3_71), .S(S_s2_80), .c_out(C_s2_80));
logic S_s2_90, C_s2_90;
FA FA_s2_90(.A(S_s3_91), .B(S_s3_90), .c_in(C_s3_81), .S(S_s2_90), .c_out(C_s2_90));
logic S_s2_100, C_s2_100;
FA FA_s2_100(.A(S_s3_101), .B(S_s3_100), .c_in(C_s3_91), .S(S_s2_100), .c_out(C_s2_100));
logic S_s2_110, C_s2_110;
FA FA_s2_110(.A(S_s3_111), .B(S_s3_110), .c_in(C_s3_101), .S(S_s2_110), .c_out(C_s2_110));
logic S_s2_120, C_s2_120;
FA FA_s2_120(.A(S_s3_121), .B(S_s3_120), .c_in(C_s3_111), .S(S_s2_120), .c_out(C_s2_120));
logic S_s2_130, C_s2_130;
FA FA_s2_130(.A(S_s3_131), .B(S_s3_130), .c_in(C_s3_121), .S(S_s2_130), .c_out(C_s2_130));
logic S_s2_140, C_s2_140;
FA FA_s2_140(.A(S_s3_141), .B(S_s3_140), .c_in(C_s3_131), .S(S_s2_140), .c_out(C_s2_140));
logic S_s2_150, C_s2_150;
FA FA_s2_150(.A(S_s3_151), .B(S_s3_150), .c_in(C_s3_141), .S(S_s2_150), .c_out(C_s2_150));
logic S_s2_160, C_s2_160;
FA FA_s2_160(.A(S_s3_161), .B(S_s3_160), .c_in(C_s3_151), .S(S_s2_160), .c_out(C_s2_160));
logic S_s2_170, C_s2_170;
FA FA_s2_170(.A(S_s3_171), .B(S_s3_170), .c_in(C_s3_161), .S(S_s2_170), .c_out(C_s2_170));
logic S_s2_180, C_s2_180;
FA FA_s2_180(.A(S_s3_181), .B(S_s3_180), .c_in(C_s3_171), .S(S_s2_180), .c_out(C_s2_180));
logic S_s2_190, C_s2_190;
FA FA_s2_190(.A(S_s3_191), .B(S_s3_190), .c_in(C_s3_181), .S(S_s2_190), .c_out(C_s2_190));
logic S_s2_200, C_s2_200;
FA FA_s2_200(.A(S_s3_201), .B(S_s3_200), .c_in(C_s3_191), .S(S_s2_200), .c_out(C_s2_200));
logic S_s2_210, C_s2_210;
FA FA_s2_210(.A(S_s3_211), .B(S_s3_210), .c_in(C_s3_201), .S(S_s2_210), .c_out(C_s2_210));
logic S_s2_220, C_s2_220;
FA FA_s2_220(.A(S_s3_221), .B(S_s3_220), .c_in(C_s3_211), .S(S_s2_220), .c_out(C_s2_220));
logic S_s2_230, C_s2_230;
FA FA_s2_230(.A(S_s3_231), .B(S_s3_230), .c_in(C_s3_221), .S(S_s2_230), .c_out(C_s2_230));
logic S_s2_240, C_s2_240;
FA FA_s2_240(.A(S_s3_241), .B(S_s3_240), .c_in(C_s3_231), .S(S_s2_240), .c_out(C_s2_240));
logic S_s2_250, C_s2_250;
FA FA_s2_250(.A(S_s3_251), .B(S_s3_250), .c_in(C_s3_241), .S(S_s2_250), .c_out(C_s2_250));
logic S_s2_260, C_s2_260;
FA FA_s2_260(.A(S_s3_261), .B(S_s3_260), .c_in(C_s3_251), .S(S_s2_260), .c_out(C_s2_260));
logic S_s2_270, C_s2_270;
FA FA_s2_270(.A(S_s3_271), .B(S_s3_270), .c_in(C_s3_261), .S(S_s2_270), .c_out(C_s2_270));
logic S_s2_280, C_s2_280;
FA FA_s2_280(.A(S_s3_281), .B(S_s3_280), .c_in(C_s3_271), .S(S_s2_280), .c_out(C_s2_280));
logic S_s2_290, C_s2_290;
FA FA_s2_290(.A(S_s3_291), .B(S_s3_290), .c_in(C_s3_281), .S(S_s2_290), .c_out(C_s2_290));
logic S_s2_300, C_s2_300;
FA FA_s2_300(.A(S_s3_301), .B(S_s3_300), .c_in(C_s3_291), .S(S_s2_300), .c_out(C_s2_300));
logic S_s2_310, C_s2_310;
FA FA_s2_310(.A(S_s3_311), .B(S_s3_310), .c_in(C_s3_301), .S(S_s2_310), .c_out(C_s2_310));
logic S_s2_320, C_s2_320;
FA FA_s2_320(.A(S_s3_321), .B(S_s3_320), .c_in(C_s3_311), .S(S_s2_320), .c_out(C_s2_320));
logic S_s2_330, C_s2_330;
FA FA_s2_330(.A(S_s3_331), .B(S_s3_330), .c_in(C_s3_321), .S(S_s2_330), .c_out(C_s2_330));
logic S_s2_340, C_s2_340;
FA FA_s2_340(.A(S_s3_341), .B(S_s3_340), .c_in(C_s3_331), .S(S_s2_340), .c_out(C_s2_340));
logic S_s2_350, C_s2_350;
FA FA_s2_350(.A(S_s3_351), .B(S_s3_350), .c_in(C_s3_341), .S(S_s2_350), .c_out(C_s2_350));
logic S_s2_360, C_s2_360;
FA FA_s2_360(.A(S_s3_361), .B(S_s3_360), .c_in(C_s3_351), .S(S_s2_360), .c_out(C_s2_360));
logic S_s2_370, C_s2_370;
FA FA_s2_370(.A(S_s3_371), .B(S_s3_370), .c_in(C_s3_361), .S(S_s2_370), .c_out(C_s2_370));
logic S_s2_380, C_s2_380;
FA FA_s2_380(.A(S_s3_381), .B(S_s3_380), .c_in(C_s3_371), .S(S_s2_380), .c_out(C_s2_380));
logic S_s2_390, C_s2_390;
FA FA_s2_390(.A(S_s3_391), .B(S_s3_390), .c_in(C_s3_381), .S(S_s2_390), .c_out(C_s2_390));
logic S_s2_400, C_s2_400;
FA FA_s2_400(.A(S_s3_401), .B(S_s3_400), .c_in(C_s3_391), .S(S_s2_400), .c_out(C_s2_400));
logic S_s2_410, C_s2_410;
FA FA_s2_410(.A(S_s3_411), .B(S_s3_410), .c_in(C_s3_401), .S(S_s2_410), .c_out(C_s2_410));
logic S_s2_420, C_s2_420;
FA FA_s2_420(.A(S_s3_421), .B(S_s3_420), .c_in(C_s3_411), .S(S_s2_420), .c_out(C_s2_420));
logic S_s2_430, C_s2_430;
FA FA_s2_430(.A(S_s3_431), .B(S_s3_430), .c_in(C_s3_421), .S(S_s2_430), .c_out(C_s2_430));
logic S_s2_440, C_s2_440;
FA FA_s2_440(.A(S_s3_441), .B(S_s3_440), .c_in(C_s3_431), .S(S_s2_440), .c_out(C_s2_440));
logic S_s2_450, C_s2_450;
FA FA_s2_450(.A(S_s3_451), .B(S_s3_450), .c_in(C_s3_441), .S(S_s2_450), .c_out(C_s2_450));
logic S_s2_460, C_s2_460;
FA FA_s2_460(.A(S_s3_461), .B(S_s3_460), .c_in(C_s3_451), .S(S_s2_460), .c_out(C_s2_460));
logic S_s2_470, C_s2_470;
FA FA_s2_470(.A(S_s3_471), .B(S_s3_470), .c_in(C_s3_461), .S(S_s2_470), .c_out(C_s2_470));
logic S_s2_480, C_s2_480;
FA FA_s2_480(.A(S_s3_481), .B(S_s3_480), .c_in(C_s3_471), .S(S_s2_480), .c_out(C_s2_480));
logic S_s2_490, C_s2_490;
FA FA_s2_490(.A(S_s3_491), .B(S_s3_490), .c_in(C_s3_481), .S(S_s2_490), .c_out(C_s2_490));
logic S_s2_500, C_s2_500;
FA FA_s2_500(.A(S_s3_501), .B(S_s3_500), .c_in(C_s3_491), .S(S_s2_500), .c_out(C_s2_500));
logic S_s2_510, C_s2_510;
FA FA_s2_510(.A(S_s3_511), .B(S_s3_510), .c_in(C_s3_501), .S(S_s2_510), .c_out(C_s2_510));
logic S_s2_520, C_s2_520;
FA FA_s2_520(.A(S_s3_521), .B(S_s3_520), .c_in(C_s3_511), .S(S_s2_520), .c_out(C_s2_520));
logic S_s2_530, C_s2_530;
FA FA_s2_530(.A(S_s3_531), .B(S_s3_530), .c_in(C_s3_521), .S(S_s2_530), .c_out(C_s2_530));
logic S_s2_540, C_s2_540;
FA FA_s2_540(.A(S_s3_541), .B(S_s3_540), .c_in(C_s3_531), .S(S_s2_540), .c_out(C_s2_540));
logic S_s2_550, C_s2_550;
FA FA_s2_550(.A(S_s3_551), .B(S_s3_550), .c_in(C_s3_541), .S(S_s2_550), .c_out(C_s2_550));
logic S_s2_560, C_s2_560;
FA FA_s2_560(.A(S_s3_561), .B(S_s3_560), .c_in(C_s3_551), .S(S_s2_560), .c_out(C_s2_560));
logic S_s2_570, C_s2_570;
FA FA_s2_570(.A(S_s3_571), .B(S_s3_570), .c_in(C_s3_561), .S(S_s2_570), .c_out(C_s2_570));
logic S_s2_580, C_s2_580;
FA FA_s2_580(.A(S_s3_581), .B(S_s3_580), .c_in(C_s3_571), .S(S_s2_580), .c_out(C_s2_580));
logic S_s2_590, C_s2_590;
FA FA_s2_590(.A(S_s3_590), .B(C_s3_581), .c_in(C_s3_580), .S(S_s2_590), .c_out(C_s2_590));
logic S_s2_600, C_s2_600;
FA FA_s2_600(.A(C_s3_590), .B(comb[29][31]), .c_in(comb[30][30]), .S(S_s2_600), .c_out(C_s2_600));
// stage 2 end ======================================================================================================= 

// stage 1 begin ======================================================================================================= 
logic S_s1_20, C_s1_20;
HA HA_s1_20(.A(comb[0][2]), .B(comb[1][1]), .S(S_s1_20), .c_out(C_s1_20));
logic S_s1_30, C_s1_30;
FA FA_s1_30(.A(S_s2_30), .B(comb[2][1]), .c_in(comb[3][0]), .S(S_s1_30), .c_out(C_s1_30));
logic S_s1_40, C_s1_40;
FA FA_s1_40(.A(S_s2_40), .B(C_s2_30), .c_in(comb[4][0]), .S(S_s1_40), .c_out(C_s1_40));
logic S_s1_50, C_s1_50;
FA FA_s1_50(.A(S_s2_50), .B(C_s2_40), .c_in(comb[5][0]), .S(S_s1_50), .c_out(C_s1_50));
logic S_s1_60, C_s1_60;
FA FA_s1_60(.A(S_s2_60), .B(C_s2_50), .c_in(C_s3_50), .S(S_s1_60), .c_out(C_s1_60));
logic S_s1_70, C_s1_70;
FA FA_s1_70(.A(S_s2_70), .B(C_s2_60), .c_in(C_s3_60), .S(S_s1_70), .c_out(C_s1_70));
logic S_s1_80, C_s1_80;
FA FA_s1_80(.A(S_s2_80), .B(C_s2_70), .c_in(C_s3_70), .S(S_s1_80), .c_out(C_s1_80));
logic S_s1_90, C_s1_90;
FA FA_s1_90(.A(S_s2_90), .B(C_s2_80), .c_in(C_s3_80), .S(S_s1_90), .c_out(C_s1_90));
logic S_s1_100, C_s1_100;
FA FA_s1_100(.A(S_s2_100), .B(C_s2_90), .c_in(C_s3_90), .S(S_s1_100), .c_out(C_s1_100));
logic S_s1_110, C_s1_110;
FA FA_s1_110(.A(S_s2_110), .B(C_s2_100), .c_in(C_s3_100), .S(S_s1_110), .c_out(C_s1_110));
logic S_s1_120, C_s1_120;
FA FA_s1_120(.A(S_s2_120), .B(C_s2_110), .c_in(C_s3_110), .S(S_s1_120), .c_out(C_s1_120));
logic S_s1_130, C_s1_130;
FA FA_s1_130(.A(S_s2_130), .B(C_s2_120), .c_in(C_s3_120), .S(S_s1_130), .c_out(C_s1_130));
logic S_s1_140, C_s1_140;
FA FA_s1_140(.A(S_s2_140), .B(C_s2_130), .c_in(C_s3_130), .S(S_s1_140), .c_out(C_s1_140));
logic S_s1_150, C_s1_150;
FA FA_s1_150(.A(S_s2_150), .B(C_s2_140), .c_in(C_s3_140), .S(S_s1_150), .c_out(C_s1_150));
logic S_s1_160, C_s1_160;
FA FA_s1_160(.A(S_s2_160), .B(C_s2_150), .c_in(C_s3_150), .S(S_s1_160), .c_out(C_s1_160));
logic S_s1_170, C_s1_170;
FA FA_s1_170(.A(S_s2_170), .B(C_s2_160), .c_in(C_s3_160), .S(S_s1_170), .c_out(C_s1_170));
logic S_s1_180, C_s1_180;
FA FA_s1_180(.A(S_s2_180), .B(C_s2_170), .c_in(C_s3_170), .S(S_s1_180), .c_out(C_s1_180));
logic S_s1_190, C_s1_190;
FA FA_s1_190(.A(S_s2_190), .B(C_s2_180), .c_in(C_s3_180), .S(S_s1_190), .c_out(C_s1_190));
logic S_s1_200, C_s1_200;
FA FA_s1_200(.A(S_s2_200), .B(C_s2_190), .c_in(C_s3_190), .S(S_s1_200), .c_out(C_s1_200));
logic S_s1_210, C_s1_210;
FA FA_s1_210(.A(S_s2_210), .B(C_s2_200), .c_in(C_s3_200), .S(S_s1_210), .c_out(C_s1_210));
logic S_s1_220, C_s1_220;
FA FA_s1_220(.A(S_s2_220), .B(C_s2_210), .c_in(C_s3_210), .S(S_s1_220), .c_out(C_s1_220));
logic S_s1_230, C_s1_230;
FA FA_s1_230(.A(S_s2_230), .B(C_s2_220), .c_in(C_s3_220), .S(S_s1_230), .c_out(C_s1_230));
logic S_s1_240, C_s1_240;
FA FA_s1_240(.A(S_s2_240), .B(C_s2_230), .c_in(C_s3_230), .S(S_s1_240), .c_out(C_s1_240));
logic S_s1_250, C_s1_250;
FA FA_s1_250(.A(S_s2_250), .B(C_s2_240), .c_in(C_s3_240), .S(S_s1_250), .c_out(C_s1_250));
logic S_s1_260, C_s1_260;
FA FA_s1_260(.A(S_s2_260), .B(C_s2_250), .c_in(C_s3_250), .S(S_s1_260), .c_out(C_s1_260));
logic S_s1_270, C_s1_270;
FA FA_s1_270(.A(S_s2_270), .B(C_s2_260), .c_in(C_s3_260), .S(S_s1_270), .c_out(C_s1_270));
logic S_s1_280, C_s1_280;
FA FA_s1_280(.A(S_s2_280), .B(C_s2_270), .c_in(C_s3_270), .S(S_s1_280), .c_out(C_s1_280));
logic S_s1_290, C_s1_290;
FA FA_s1_290(.A(S_s2_290), .B(C_s2_280), .c_in(C_s3_280), .S(S_s1_290), .c_out(C_s1_290));
logic S_s1_300, C_s1_300;
FA FA_s1_300(.A(S_s2_300), .B(C_s2_290), .c_in(C_s3_290), .S(S_s1_300), .c_out(C_s1_300));
logic S_s1_310, C_s1_310;
FA FA_s1_310(.A(S_s2_310), .B(C_s2_300), .c_in(C_s3_300), .S(S_s1_310), .c_out(C_s1_310));
logic S_s1_320, C_s1_320;
FA FA_s1_320(.A(S_s2_320), .B(C_s2_310), .c_in(C_s3_310), .S(S_s1_320), .c_out(C_s1_320));
logic S_s1_330, C_s1_330;
FA FA_s1_330(.A(S_s2_330), .B(C_s2_320), .c_in(C_s3_320), .S(S_s1_330), .c_out(C_s1_330));
logic S_s1_340, C_s1_340;
FA FA_s1_340(.A(S_s2_340), .B(C_s2_330), .c_in(C_s3_330), .S(S_s1_340), .c_out(C_s1_340));
logic S_s1_350, C_s1_350;
FA FA_s1_350(.A(S_s2_350), .B(C_s2_340), .c_in(C_s3_340), .S(S_s1_350), .c_out(C_s1_350));
logic S_s1_360, C_s1_360;
FA FA_s1_360(.A(S_s2_360), .B(C_s2_350), .c_in(C_s3_350), .S(S_s1_360), .c_out(C_s1_360));
logic S_s1_370, C_s1_370;
FA FA_s1_370(.A(S_s2_370), .B(C_s2_360), .c_in(C_s3_360), .S(S_s1_370), .c_out(C_s1_370));
logic S_s1_380, C_s1_380;
FA FA_s1_380(.A(S_s2_380), .B(C_s2_370), .c_in(C_s3_370), .S(S_s1_380), .c_out(C_s1_380));
logic S_s1_390, C_s1_390;
FA FA_s1_390(.A(S_s2_390), .B(C_s2_380), .c_in(C_s3_380), .S(S_s1_390), .c_out(C_s1_390));
logic S_s1_400, C_s1_400;
FA FA_s1_400(.A(S_s2_400), .B(C_s2_390), .c_in(C_s3_390), .S(S_s1_400), .c_out(C_s1_400));
logic S_s1_410, C_s1_410;
FA FA_s1_410(.A(S_s2_410), .B(C_s2_400), .c_in(C_s3_400), .S(S_s1_410), .c_out(C_s1_410));
logic S_s1_420, C_s1_420;
FA FA_s1_420(.A(S_s2_420), .B(C_s2_410), .c_in(C_s3_410), .S(S_s1_420), .c_out(C_s1_420));
logic S_s1_430, C_s1_430;
FA FA_s1_430(.A(S_s2_430), .B(C_s2_420), .c_in(C_s3_420), .S(S_s1_430), .c_out(C_s1_430));
logic S_s1_440, C_s1_440;
FA FA_s1_440(.A(S_s2_440), .B(C_s2_430), .c_in(C_s3_430), .S(S_s1_440), .c_out(C_s1_440));
logic S_s1_450, C_s1_450;
FA FA_s1_450(.A(S_s2_450), .B(C_s2_440), .c_in(C_s3_440), .S(S_s1_450), .c_out(C_s1_450));
logic S_s1_460, C_s1_460;
FA FA_s1_460(.A(S_s2_460), .B(C_s2_450), .c_in(C_s3_450), .S(S_s1_460), .c_out(C_s1_460));
logic S_s1_470, C_s1_470;
FA FA_s1_470(.A(S_s2_470), .B(C_s2_460), .c_in(C_s3_460), .S(S_s1_470), .c_out(C_s1_470));
logic S_s1_480, C_s1_480;
FA FA_s1_480(.A(S_s2_480), .B(C_s2_470), .c_in(C_s3_470), .S(S_s1_480), .c_out(C_s1_480));
logic S_s1_490, C_s1_490;
FA FA_s1_490(.A(S_s2_490), .B(C_s2_480), .c_in(C_s3_480), .S(S_s1_490), .c_out(C_s1_490));
logic S_s1_500, C_s1_500;
FA FA_s1_500(.A(S_s2_500), .B(C_s2_490), .c_in(C_s3_490), .S(S_s1_500), .c_out(C_s1_500));
logic S_s1_510, C_s1_510;
FA FA_s1_510(.A(S_s2_510), .B(C_s2_500), .c_in(C_s3_500), .S(S_s1_510), .c_out(C_s1_510));
logic S_s1_520, C_s1_520;
FA FA_s1_520(.A(S_s2_520), .B(C_s2_510), .c_in(C_s3_510), .S(S_s1_520), .c_out(C_s1_520));
logic S_s1_530, C_s1_530;
FA FA_s1_530(.A(S_s2_530), .B(C_s2_520), .c_in(C_s3_520), .S(S_s1_530), .c_out(C_s1_530));
logic S_s1_540, C_s1_540;
FA FA_s1_540(.A(S_s2_540), .B(C_s2_530), .c_in(C_s3_530), .S(S_s1_540), .c_out(C_s1_540));
logic S_s1_550, C_s1_550;
FA FA_s1_550(.A(S_s2_550), .B(C_s2_540), .c_in(C_s3_540), .S(S_s1_550), .c_out(C_s1_550));
logic S_s1_560, C_s1_560;
FA FA_s1_560(.A(S_s2_560), .B(C_s2_550), .c_in(C_s3_550), .S(S_s1_560), .c_out(C_s1_560));
logic S_s1_570, C_s1_570;
FA FA_s1_570(.A(S_s2_570), .B(C_s2_560), .c_in(C_s3_560), .S(S_s1_570), .c_out(C_s1_570));
logic S_s1_580, C_s1_580;
FA FA_s1_580(.A(S_s2_580), .B(C_s2_570), .c_in(C_s3_570), .S(S_s1_580), .c_out(C_s1_580));
logic S_s1_590, C_s1_590;
FA FA_s1_590(.A(S_s2_590), .B(C_s2_580), .c_in(comb[31][28]), .S(S_s1_590), .c_out(C_s1_590));
logic S_s1_600, C_s1_600;
FA FA_s1_600(.A(S_s2_600), .B(C_s2_590), .c_in(comb[31][29]), .S(S_s1_600), .c_out(C_s1_600));
logic S_s1_610, C_s1_610;
FA FA_s1_610(.A(C_s2_600), .B(comb[30][31]), .c_in(comb[31][30]), .S(S_s1_610), .c_out(C_s1_610));
// stage 1 end ======================================================================================================= 


logic [63:0] last_top_row, last_bot_row;
assign last_top_row = {1'b0, C_s1_610, S_s1_610, S_s1_600, S_s1_590, S_s1_580, S_s1_570, S_s1_560, S_s1_550, S_s1_540, S_s1_530, S_s1_520, S_s1_510, S_s1_500, S_s1_490, S_s1_480, S_s1_470, S_s1_460, S_s1_450, S_s1_440, S_s1_430, S_s1_420, S_s1_410, S_s1_400, S_s1_390, S_s1_380, S_s1_370, S_s1_360, S_s1_350, S_s1_340, S_s1_330, S_s1_320, S_s1_310, S_s1_300, S_s1_290, S_s1_280, S_s1_270, S_s1_260, S_s1_250, S_s1_240, S_s1_230, S_s1_220, S_s1_210, S_s1_200, S_s1_190, S_s1_180, S_s1_170, S_s1_160, S_s1_150, S_s1_140, S_s1_130, S_s1_120, S_s1_110, S_s1_100, S_s1_90, S_s1_80, S_s1_70, S_s1_60, S_s1_50, S_s1_40, S_s1_30, S_s1_20, comb[0][1], comb[0][0]};
assign last_bot_row = {1'b0, comb[31][31], C_s1_600, C_s1_590, C_s1_580, C_s1_570, C_s1_560, C_s1_550, C_s1_540, C_s1_530, C_s1_520, C_s1_510, C_s1_500, C_s1_490, C_s1_480, C_s1_470, C_s1_460, C_s1_450, C_s1_440, C_s1_430, C_s1_420, C_s1_410, C_s1_400, C_s1_390, C_s1_380, C_s1_370, C_s1_360, C_s1_350, C_s1_340, C_s1_330, C_s1_320, C_s1_310, C_s1_300, C_s1_290, C_s1_280, C_s1_270, C_s1_260, C_s1_250, C_s1_240, C_s1_230, C_s1_220, C_s1_210, C_s1_200, C_s1_190, C_s1_180, C_s1_170, C_s1_160, C_s1_150, C_s1_140, C_s1_130, C_s1_120, C_s1_110, C_s1_100, C_s1_90, C_s1_80, C_s1_70, C_s1_60, C_s1_50, C_s1_40, C_s1_30, C_s1_20, comb[2][0], comb[1][0], 1'b0};
assign prodAB = last_top_row + last_bot_row;    // combine and find the sum, naive implementation
endmodule
